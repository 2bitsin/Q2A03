
module core_decoder(I_ir, I_t, O_control);
	input wire[7:0] I_ir;
	input wire[3:0] I_t;
	output wire[92:0] O_control;
	
	wire w000 = (I_ir ==? 8'b0?101?00);
	wire w001 = (I_ir ==? 8'b0??0000?);
	wire w002 = (I_ir ==? 8'b0???0?11);
	wire w003 = (I_ir ==? 8'b0????110);
	wire w004 = (I_ir ==? 8'b1001??01);
	wire w005 = (I_ir ==? 8'b11?011??);
	wire w006 = (I_ir ==? 8'b?0?000?1);
	wire w007 = (I_ir ==? 8'b?0?011??);
	wire w008 = (I_ir ==? 8'b?0??0001);
	wire w009 = (I_ir ==? 8'b?1?011?1);
	wire w010 = (I_ir ==? 8'b?1?0?11?);
	wire w011 = (I_ir ==? 8'b?1??00?1);
	wire w012 = (I_ir ==? 8'b?1???110);
	wire w013 = (I_ir ==? 8'b??1?00?1);
	wire w014 = (I_ir ==? 8'b???101??);
	wire w015 = (I_ir ==? 8'b0??0??00);
	wire w016 = (I_ir ==? 8'b0??1???1);
	wire w017 = (I_ir ==? 8'b0????1??);
	wire w018 = (I_ir ==? 8'b101?0??1);
	wire w019 = (I_ir ==? 8'b?1?111??);
	wire w020 = (I_ir ==? 8'b?1?1???1);
	wire w021 = (I_ir ==? 8'b??1111??);
	wire w022 = (I_ir ==? 8'b???00??1);
	wire w023 = (I_ir ==? 8'b???0?1??);
	wire w024 = (I_ir ==? 8'b???1??01);
	wire w025 = (I_ir ==? 8'b????01??);
	wire w026 = (I_ir ==? 8'b011?11?0);
	wire w027 = (I_ir ==? 8'b0??111??);
	wire w028 = (I_ir ==? 8'b0??11?11);
	wire w029 = (I_ir ==? 8'b0????11?);
	wire w030 = (I_ir ==? 8'b100?0001);
	wire w031 = (I_ir ==? 8'b?1?11?11);
	wire w032 = (I_ir ==? 8'b?1???11?);
	wire w033 = (I_ir ==? 8'b???000?1);
	wire w034 = (I_ir ==? 8'b???11?01);
	wire w035 = (I_ir ==? 8'b0??1?11?);
	wire w036 = (I_ir ==? 8'b0??1??11);
	wire w037 = (I_ir ==? 8'b0???111?);
	wire w038 = (I_ir ==? 8'b101?00?1);
	wire w039 = (I_ir ==? 8'b11?1?011);
	wire w040 = (I_ir ==? 8'b?1?1?11?);
	wire w041 = (I_ir ==? 8'b?1??111?);
	wire w042 = (I_ir ==? 8'b????0001);
	wire w043 = (I_ir ==? 8'b0???0011);
	wire w044 = (I_ir ==? 8'b?1??0011);
	wire w045 = (I_ir ==? 8'b00000000);
	wire w046 = (I_ir ==? 8'b00?1111?);
	wire w047 = (I_ir ==? 8'b00??0011);
	wire w048 = (I_ir ==? 8'b?1?1111?);
	wire w049 = (I_ir ==? 8'b?1?1?011);
	wire w050 = (I_ir ==? 8'b0?101000);
	wire w051 = (I_ir ==? 8'b0??00000);
	wire w052 = (I_ir ==? 8'b0??0?000);
	wire w053 = (I_ir ==? 8'b01000000);
	wire w054 = (I_ir ==? 8'b00?00000);
	wire w055 = (I_ir ==? 8'b0??0011?);
	wire w056 = (I_ir ==? 8'b100011??);
	wire w057 = (I_ir ==? 8'b100101??);
	wire w058 = (I_ir ==? 8'b?1?0011?);
	wire w059 = (I_ir ==? 8'b0??11110);
	wire w060 = (I_ir ==? 8'b11?1111?);
	wire w061 = (I_ir ==? 8'b00?0?110);
	wire w062 = (I_ir ==? 8'b0??01111);
	wire w063 = (I_ir ==? 8'b0??1011?);
	wire w064 = (I_ir ==? 8'b10011?01);
	wire w065 = (I_ir ==? 8'b11??011?);
	wire w066 = (I_ir ==? 8'b?1?0111?);
	wire w067 = (I_ir ==? 8'b?1??0110);
	wire w068 = (I_ir ==? 8'b00?10110);
	wire w069 = (I_ir ==? 8'b0???1110);
	wire w070 = (I_ir ==? 8'b100000?1);
	wire w071 = (I_ir ==? 8'b11?1?11?);
	wire w072 = (I_ir ==? 8'b11??111?);
	wire w073 = (I_ir ==? 8'b?1?1?110);
	wire w074 = (I_ir ==? 8'b11??0011);
	wire w075 = (I_ir ==? 8'b0?001000);
	wire w076 = (I_ir ==? 8'b100001??);
	wire w077 = (I_ir ==? 8'b11001011);
	wire w078 = (I_ir ==? 8'b00100000);
	wire w079 = (I_ir ==? 8'b0000?000);
	wire w080 = (I_ir ==? 8'b00001000);
	wire w081 = (I_ir ==? 8'b00100?00);
	wire w082 = (I_ir ==? 8'b001011??);
	wire w083 = (I_ir ==? 8'b0?00?1??);
	wire w084 = (I_ir ==? 8'b0??10??1);
	wire w085 = (I_ir ==? 8'b11010??1);
	wire w086 = (I_ir ==? 8'b1??011??);
	wire w087 = (I_ir ==? 8'b?0?10001);
	wire w088 = (I_ir ==? 8'b?110?11?);
	wire w089 = (I_ir ==? 8'b??110??1);
	wire w090 = (I_ir ==? 8'b???0?1?1);
	wire w091 = (I_ir ==? 8'b01101100);
	wire w092 = (I_ir ==? 8'b00?11??1);
	wire w093 = (I_ir ==? 8'b0?0?11??);
	wire w094 = (I_ir ==? 8'b0?1?11?1);
	wire w095 = (I_ir ==? 8'b?01?11??);
	wire w096 = (I_ir ==? 8'b??1?111?);
	wire w097 = (I_ir ==? 8'b0??100?1);
	wire w098 = (I_ir ==? 8'b101100?1);
	wire w099 = (I_ir ==? 8'b?1?100?1);
	wire w100 = (I_ir ==? 8'b???10001);
	wire w101 = (I_ir ==? 8'b01001100);
	wire w102 = (I_ir ==? 8'b0010000?);
	wire w103 = (I_ir ==? 8'b01?0000?);
	wire w104 = (I_ir ==? 8'b0??0111?);
	wire w105 = (I_ir ==? 8'b10?000?1);
	wire w106 = (I_ir ==? 8'b?1?1011?);
	wire w107 = (I_ir ==? 8'b00?0110?);
	wire w108 = (I_ir ==? 8'b10?011??);
	wire w109 = (I_ir ==? 8'b10?101??);
	wire w110 = (I_ir ==? 8'b1??0110?);
	wire w111 = (I_ir ==? 8'b???01101);
	wire w112 = (I_ir ==? 8'b???1010?);
	wire w113 = (I_ir ==? 8'b???10?00);
	wire w114 = (I_ir ==? 8'b1010?0?0);
	wire w115 = (I_ir ==? 8'b10?0?000);
	wire w116 = (I_ir ==? 8'b11?010??);
	wire w117 = (I_ir ==? 8'b11?0?0?0);
	wire w118 = (I_ir ==? 8'b1?1010?1);
	wire w119 = (I_ir ==? 8'b1???10?0);
	wire w120 = (I_ir ==? 8'b???01001);
	wire w121 = (I_ir ==? 8'b???110?0);
	wire w122 = (I_ir ==? 8'b????1010);
	wire w123 = (I_ir ==? 8'b00?0011?);
	wire w124 = (I_ir ==? 8'b011?1100);
	wire w125 = (I_ir ==? 8'b0??1110?);
	wire w126 = (I_ir ==? 8'b101111??);
	wire w127 = (I_ir ==? 8'b11?1110?);
	wire w128 = (I_ir ==? 8'b0100?100);
	wire w129 = (I_ir ==? 8'b10?001??);
	wire w130 = (I_ir ==? 8'b???0010?);
	wire w131 = (I_ir ==? 8'b101010?1);
	wire w132 = (I_ir ==? 8'b11000?1?);
	wire w133 = (I_ir ==? 8'b11?0?0?1);
	wire w134 = (I_ir ==? 8'b1?10001?);
	wire w135 = (I_ir ==? 8'b1?110??1);
	wire w136 = (I_ir ==? 8'b1??0000?);
	wire w137 = (I_ir ==? 8'b1??0?1??);
	wire w138 = (I_ir ==? 8'b?01?000?);
	wire w139 = (I_ir ==? 8'b???1000?);
	wire w140 = (I_ir ==? 8'b??????01);
	wire w141 = (I_ir ==? 8'b01??11?1);
	wire w142 = (I_ir ==? 8'b0?0111??);
	wire w143 = (I_ir ==? 8'b0?0?111?);
	wire w144 = (I_ir ==? 8'b0??11??1);
	wire w145 = (I_ir ==? 8'b110?11??);
	wire w146 = (I_ir ==? 8'b11?11?11);
	wire w147 = (I_ir ==? 8'b??1?11??);
	wire w148 = (I_ir ==? 8'b01100000);
	wire w149 = (I_ir ==? 8'b?1?11??1);
	wire w150 = (I_ir ==? 8'b0???00?1);
	wire w151 = (I_ir ==? 8'b11??00?1);
	wire w152 = (I_ir ==? 8'b0??1?1??);
	wire w153 = (I_ir ==? 8'b1?11110?);
	wire w154 = (I_ir ==? 8'b1??1?101);
	wire w155 = (I_ir ==? 8'b?1?1?1??);
	wire w156 = (I_ir ==? 8'b00???11?);
	wire w157 = (I_ir ==? 8'b11??11??);
	wire w158 = (I_ir ==? 8'b1?110?11);
	wire w159 = (I_ir ==? 8'b1??1011?);
	wire w160 = (I_ir ==? 8'b??11?1??);
	wire w161 = (I_ir ==? 8'b???10?0?);
	wire w162 = (I_ir ==? 8'b???1?001);
	wire w163 = (I_ir ==? 8'b????1101);
	wire w164 = (I_ir ==? 8'b?1?1??11);
	wire w165 = (I_ir ==? 8'b??1100?1);
	wire w166 = (I_ir ==? 8'b000111??);
	wire w167 = (I_ir ==? 8'b??110011);
	wire w168 = (I_ir ==? 8'b00?11011);
	wire w169 = (I_ir ==? 8'b0??1111?);
	wire w170 = (I_ir ==? 8'b0?010?11);
	wire w171 = (I_ir ==? 8'b?0110?11);
	wire w172 = (I_ir ==? 8'b?1?10?11);
	wire w173 = (I_ir ==? 8'b00001111);
	wire w174 = (I_ir ==? 8'b00010111);
	wire w175 = (I_ir ==? 8'b000?0001);
	wire w176 = (I_ir ==? 8'b00011?11);
	wire w177 = (I_ir ==? 8'b000?0011);
	wire w178 = (I_ir ==? 8'b00000111);
	wire w179 = (I_ir ==? 8'b00011?01);
	wire w180 = (I_ir ==? 8'b00001001);
	wire w181 = (I_ir ==? 8'b00001101);
	wire w182 = (I_ir ==? 8'b00010101);
	wire w183 = (I_ir ==? 8'b00000101);
	wire w184 = (I_ir ==? 8'b001?0001);
	wire w185 = (I_ir ==? 8'b0??10111);
	wire w186 = (I_ir ==? 8'b?11?0001);
	wire w187 = (I_ir ==? 8'b??0?0001);
	wire w188 = (I_ir ==? 8'b0010110?);
	wire w189 = (I_ir ==? 8'b00?01101);
	wire w190 = (I_ir ==? 8'b0??10101);
	wire w191 = (I_ir ==? 8'b100011?1);
	wire w192 = (I_ir ==? 8'b100101?1);
	wire w193 = (I_ir ==? 8'b11?00111);
	wire w194 = (I_ir ==? 8'b?1?01101);
	wire w195 = (I_ir ==? 8'b?1?10101);
	wire w196 = (I_ir ==? 8'b??010101);
	wire w197 = (I_ir ==? 8'b00111?01);
	wire w198 = (I_ir ==? 8'b0??00111);
	wire w199 = (I_ir ==? 8'b11?01111);
	wire w200 = (I_ir ==? 8'b11?10111);
	wire w201 = (I_ir ==? 8'b?1?11?01);
	wire w202 = (I_ir ==? 8'b??011?01);
	wire w203 = (I_ir ==? 8'b0??01001);
	wire w204 = (I_ir ==? 8'b0??01010);
	wire w205 = (I_ir ==? 8'b101010?0);
	wire w206 = (I_ir ==? 8'b11?010?1);
	wire w207 = (I_ir ==? 8'b0010010?);
	wire w208 = (I_ir ==? 8'b01001000);
	wire w209 = (I_ir ==? 8'b0??00101);
	wire w210 = (I_ir ==? 8'b100001?1);
	wire w211 = (I_ir ==? 8'b11?00101);
	wire w212 = (I_ir ==? 8'b?1??0001);
	wire w213 = (I_ir ==? 8'b??1?0001);
	wire w214 = (I_ir ==? 8'b00?10101);
	wire w215 = (I_ir ==? 8'b01101000);
	wire w216 = (I_ir ==? 8'b0??01101);
	wire w217 = (I_ir ==? 8'b101011??);
	wire w218 = (I_ir ==? 8'b101101??);
	wire w219 = (I_ir ==? 8'b11?0110?);
	wire w220 = (I_ir ==? 8'b0??11?01);
	wire w221 = (I_ir ==? 8'b1?111?01);
	wire w222 = (I_ir ==? 8'b101000?0);
	wire w223 = (I_ir ==? 8'b11?00000);
	wire w224 = (I_ir ==? 8'b1?100000);
	wire w225 = (I_ir ==? 8'b?1?01001);
	wire w226 = (I_ir ==? 8'b101001??);
	wire w227 = (I_ir ==? 8'b11?0010?);
	wire w228 = (I_ir ==? 8'b?010010?);
	wire w229 = (I_ir ==? 8'b?1?00101);
	wire w230 = (I_ir ==? 8'b0???0001);
	wire w231 = (I_ir ==? 8'b11111?11);
	wire w232 = (I_ir ==? 8'b101011?1);
	wire w233 = (I_ir ==? 8'b101101?1);
	wire w234 = (I_ir ==? 8'b11100111);
	wire w235 = (I_ir ==? 8'b1?101101);
	wire w236 = (I_ir ==? 8'b??110101);
	wire w237 = (I_ir ==? 8'b101111?1);
	wire w238 = (I_ir ==? 8'b11101111);
	wire w239 = (I_ir ==? 8'b11110111);
	wire w240 = (I_ir ==? 8'b??111?01);
	wire w241 = (I_ir ==? 8'b111?0011);
	wire w242 = (I_ir ==? 8'b10011000);
	wire w243 = (I_ir ==? 8'b?0001010);
	wire w244 = (I_ir ==? 8'b101001?1);
	wire w245 = (I_ir ==? 8'b1?100101);
	wire w246 = (I_ir ==? 8'b00000110);
	wire w247 = (I_ir ==? 8'b0000?110);
	wire w248 = (I_ir ==? 8'b000?0110);
	wire w249 = (I_ir ==? 8'b0001?110);
	wire w250 = (I_ir ==? 8'b000?1110);
	wire w251 = (I_ir ==? 8'b00001010);
	wire w252 = (I_ir ==? 8'b00011110);
	wire w253 = (I_ir ==? 8'b00?10111);
	wire w254 = (I_ir ==? 8'b?1?01111);
	wire w255 = (I_ir ==? 8'b?1?10111);
	wire w256 = (I_ir ==? 8'b0?100110);
	wire w257 = (I_ir ==? 8'b11?00110);
	wire w258 = (I_ir ==? 8'b?1100110);
	wire w259 = (I_ir ==? 8'b0?111110);
	wire w260 = (I_ir ==? 8'b11?11110);
	wire w261 = (I_ir ==? 8'b?1111110);
	wire w262 = (I_ir ==? 8'b0?101110);
	wire w263 = (I_ir ==? 8'b0?110110);
	wire w264 = (I_ir ==? 8'b11?01110);
	wire w265 = (I_ir ==? 8'b11?10110);
	wire w266 = (I_ir ==? 8'b?1101110);
	wire w267 = (I_ir ==? 8'b?1110110);
	wire w268 = (I_ir ==? 8'b0?10011?);
	wire w269 = (I_ir ==? 8'b11?0011?);
	wire w270 = (I_ir ==? 8'b?1?00111);
	wire w271 = (I_ir ==? 8'b0?001111);
	wire w272 = (I_ir ==? 8'b0?10111?);
	wire w273 = (I_ir ==? 8'b0?11011?);
	wire w274 = (I_ir ==? 8'b0?1?0110);
	wire w275 = (I_ir ==? 8'b11?0?11?);
	wire w276 = (I_ir ==? 8'b11?1011?);
	wire w277 = (I_ir ==? 8'b0?11?110);
	wire w278 = (I_ir ==? 8'b0?1?1110);
	wire w279 = (I_ir ==? 8'b00?10??1);
	wire w280 = (I_ir ==? 8'b1??10001);
	wire w281 = (I_ir ==? 8'b?1010??1);
	wire w282 = (I_ir ==? 8'b0??01110);
	wire w283 = (I_ir ==? 8'b?1?01110);
	wire w284 = (I_ir ==? 8'b?1?10110);
	wire w285 = (I_ir ==? 8'b0??00110);
	wire w286 = (I_ir ==? 8'b00111110);
	wire w287 = (I_ir ==? 8'b0?01?110);
	wire w288 = (I_ir ==? 8'b0?0?1110);
	wire w289 = (I_ir ==? 8'b?1?11110);
	wire w290 = (I_ir ==? 8'b0?00?110);
	wire w291 = (I_ir ==? 8'b0??10110);
	wire w292 = (I_ir ==? 8'b0?011110);
	wire w293 = (I_ir ==? 8'b0?000110);
	wire w294 = (I_ir ==? 8'b0?001110);
	wire w295 = (I_ir ==? 8'b0?0?0110);
	wire w296 = (I_ir ==? 8'b00010000);
	wire w297 = (I_ir ==? 8'b???10000);
	wire w298 = (I_ir ==? 8'b1?11?1??);
	wire w299 = (I_ir ==? 8'b11?10??1);
	wire w300 = (I_ir ==? 8'b???10?01);
	wire w301 = (I_ir ==? 8'b0??110?1);
	wire w302 = (I_ir ==? 8'b1011?11?);
	wire w303 = (I_ir ==? 8'b10?1011?);
	wire w304 = (I_ir ==? 8'b?1?110?1);
	wire w305 = (I_ir ==? 8'b???11001);
	wire w306 = (I_ir ==? 8'b0?01110?);
	wire w307 = (I_ir ==? 8'b?101110?);
	wire w308 = (I_ir ==? 8'b??11110?);
	wire w309 = (I_ir ==? 8'b00011000);
	wire w310 = (I_ir ==? 8'b00100111);
	wire w311 = (I_ir ==? 8'b00101111);
	wire w312 = (I_ir ==? 8'b00110111);
	wire w313 = (I_ir ==? 8'b10000011);
	wire w314 = (I_ir ==? 8'b001?0011);
	wire w315 = (I_ir ==? 8'b00101101);
	wire w316 = (I_ir ==? 8'b00110101);
	wire w317 = (I_ir ==? 8'b10001111);
	wire w318 = (I_ir ==? 8'b10010111);
	wire w319 = (I_ir ==? 8'b00101001);
	wire w320 = (I_ir ==? 8'b00111?11);
	wire w321 = (I_ir ==? 8'b00100101);
	wire w322 = (I_ir ==? 8'b10000111);
	wire w323 = (I_ir ==? 8'b00101110);
	wire w324 = (I_ir ==? 8'b00110110);
	wire w325 = (I_ir ==? 8'b00100110);
	wire w326 = (I_ir ==? 8'b00101010);
	wire w327 = (I_ir ==? 8'b00100100);
	wire w328 = (I_ir ==? 8'b00101100);
	wire w329 = (I_ir ==? 8'b01?00000);
	wire w330 = (I_ir ==? 8'b00101000);
	wire w331 = (I_ir ==? 8'b00110000);
	wire w332 = (I_ir ==? 8'b00111000);
	wire w333 = (I_ir ==? 8'b01001111);
	wire w334 = (I_ir ==? 8'b01010111);
	wire w335 = (I_ir ==? 8'b010?0001);
	wire w336 = (I_ir ==? 8'b01001001);
	wire w337 = (I_ir ==? 8'b01000111);
	wire w338 = (I_ir ==? 8'b01011?01);
	wire w339 = (I_ir ==? 8'b01001101);
	wire w340 = (I_ir ==? 8'b01010101);
	wire w341 = (I_ir ==? 8'b010?0011);
	wire w342 = (I_ir ==? 8'b01000101);
	wire w343 = (I_ir ==? 8'b01011?11);
	wire w344 = (I_ir ==? 8'b01000110);
	wire w345 = (I_ir ==? 8'b0101?110);
	wire w346 = (I_ir ==? 8'b010?1110);
	wire w347 = (I_ir ==? 8'b0100?110);
	wire w348 = (I_ir ==? 8'b010?0110);
	wire w349 = (I_ir ==? 8'b01001010);
	wire w350 = (I_ir ==? 8'b01011110);
	wire w351 = (I_ir ==? 8'b01010000);
	wire w352 = (I_ir ==? 8'b01011000);
	wire w353 = (I_ir ==? 8'b01101101);
	wire w354 = (I_ir ==? 8'b01110101);
	wire w355 = (I_ir ==? 8'b01101111);
	wire w356 = (I_ir ==? 8'b01110111);
	wire w357 = (I_ir ==? 8'b011?0001);
	wire w358 = (I_ir ==? 8'b01100101);
	wire w359 = (I_ir ==? 8'b01100111);
	wire w360 = (I_ir ==? 8'b01111?01);
	wire w361 = (I_ir ==? 8'b01111?11);
	wire w362 = (I_ir ==? 8'b011?0011);
	wire w363 = (I_ir ==? 8'b01101001);
	wire w364 = (I_ir ==? 8'b01100110);
	wire w365 = (I_ir ==? 8'b01101110);
	wire w366 = (I_ir ==? 8'b01110110);
	wire w367 = (I_ir ==? 8'b01101010);
	wire w368 = (I_ir ==? 8'b01111110);
	wire w369 = (I_ir ==? 8'b10111?01);
	wire w370 = (I_ir ==? 8'b01110000);
	wire w371 = (I_ir ==? 8'b01111000);
	wire w372 = (I_ir ==? 8'b10010100);
	wire w373 = (I_ir ==? 8'b1?001100);
	wire w374 = (I_ir ==? 8'b100?1000);
	wire w375 = (I_ir ==? 8'b1100?000);
	wire w376 = (I_ir ==? 8'b1?001000);
	wire w377 = (I_ir ==? 8'b1?000100);
	wire w378 = (I_ir ==? 8'b10000110);
	wire w379 = (I_ir ==? 8'b11100100);
	wire w380 = (I_ir ==? 8'b10001110);
	wire w381 = (I_ir ==? 8'b10010110);
	wire w382 = (I_ir ==? 8'b11101100);
	wire w383 = (I_ir ==? 8'b1110?000);
	wire w384 = (I_ir ==? 8'b1?001010);
	wire w385 = (I_ir ==? 8'b11011110);
	wire w386 = (I_ir ==? 8'b110?0011);
	wire w387 = (I_ir ==? 8'b11000111);
	wire w388 = (I_ir ==? 8'b11001110);
	wire w389 = (I_ir ==? 8'b11010110);
	wire w390 = (I_ir ==? 8'b11011?11);
	wire w391 = (I_ir ==? 8'b11000110);
	wire w392 = (I_ir ==? 8'b11001111);
	wire w393 = (I_ir ==? 8'b11010111);
	wire w394 = (I_ir ==? 8'b10001000);
	wire w395 = (I_ir ==? 8'b11001010);
	wire w396 = (I_ir ==? 8'b10100100);
	wire w397 = (I_ir ==? 8'b1010?000);
	wire w398 = (I_ir ==? 8'b10101100);
	wire w399 = (I_ir ==? 8'b10110100);
	wire w400 = (I_ir ==? 8'b10111100);
	wire w401 = (I_ir ==? 8'b101?1010);
	wire w402 = (I_ir ==? 8'b10?01010);
	wire w403 = (I_ir ==? 8'b10010000);
	wire w404 = (I_ir ==? 8'b10011010);
	wire w405 = (I_ir ==? 8'b1010101?);
	wire w406 = (I_ir ==? 8'b1010?010);
	wire w407 = (I_ir ==? 8'b11101000);
	wire w408 = (I_ir ==? 8'b1010111?);
	wire w409 = (I_ir ==? 8'b1011011?);
	wire w410 = (I_ir ==? 8'b1011111?);
	wire w411 = (I_ir ==? 8'b1010011?);
	wire w412 = (I_ir ==? 8'b101?0011);
	wire w413 = (I_ir ==? 8'b10110000);
	wire w414 = (I_ir ==? 8'b10111000);
	wire w415 = (I_ir ==? 8'b10111010);
	wire w416 = (I_ir ==? 8'b1100010?);
	wire w417 = (I_ir ==? 8'b11?00100);
	wire w418 = (I_ir ==? 8'b1100110?);
	wire w419 = (I_ir ==? 8'b11010101);
	wire w420 = (I_ir ==? 8'b11?01100);
	wire w421 = (I_ir ==? 8'b11011?01);
	wire w422 = (I_ir ==? 8'b11001001);
	wire w423 = (I_ir ==? 8'b110?0001);
	wire w424 = (I_ir ==? 8'b11101110);
	wire w425 = (I_ir ==? 8'b11110110);
	wire w426 = (I_ir ==? 8'b11100110);
	wire w427 = (I_ir ==? 8'b11111110);
	wire w428 = (I_ir ==? 8'b11?01000);
	wire w429 = (I_ir ==? 8'b11010000);
	wire w430 = (I_ir ==? 8'b11011000);
	wire w431 = (I_ir ==? 8'b11101101);
	wire w432 = (I_ir ==? 8'b11110101);
	wire w433 = (I_ir ==? 8'b111?0001);
	wire w434 = (I_ir ==? 8'b11111?01);
	wire w435 = (I_ir ==? 8'b111010?1);
	wire w436 = (I_ir ==? 8'b11100101);
	wire w437 = (I_ir ==? 8'b11110000);
	wire w438 = (I_ir ==? 8'b11111000);
	
	wire t0 = (I_t == 4'd0);
	wire t1 = (I_t == 4'd1);
	wire t2 = (I_t == 4'd2);
	wire t3 = (I_t == 4'd3);
	wire t4 = (I_t == 4'd4);
	wire t5 = (I_t == 4'd5);
	wire t6 = (I_t == 4'd6);
	wire t7 = (I_t == 4'd7);
	
	wire x000 = w000|w001|w002|w003|w004|w005|w006|w007|w008|w009|w010|w011|w012|w013|w014;
	wire x001 = w015|w016|w017|w018|w019|w020|w021|w022|w023|w024|w025;
	wire x002 = w026|w001|w027|w028|w029|w030|w019|w031|w032|w021|w033|w034;
	wire x003 = w001|w035|w036|w037|w038|w039|w040|w041|w033|w042;
	wire x004 = w043|w044;
	wire x005 = w045|w046|w047|w028|w048|w049|w044;
	wire x006 = w050|w051;
	wire x007 = w052;
	wire x008 = w051;
	wire x009 = w053;
	wire x010 = w054|w055|w056|w057|w058;
	wire x011 = w047|w059|w060|w039|w044;
	wire x012 = w054|w061|w062|w063|w064|w065|w066|w067;
	wire x013 = w068|w028|w069|w070|w030|w071|w072|w031|w073;
	wire x014 = w074;
	wire x015 = w045|w075|w076;
	wire x016 = w077;
	wire x017 = w045;
	wire x018 = w078;
	wire x019 = w079|w075;
	wire x020 = w054;
	wire x021 = w080;
	wire x022 = w081|w082|w083|w084|w085|w086|w087|w088|w089|w090|w025;
	wire x023 = w091|w033;
	wire x024 = w092|w093|w094|w086|w095|w019|w031|w096|w034;
	wire x025 = w097|w098|w099|w100;
	wire x026 = w101;
	wire x027 = w091;
	wire x028 = w102|w103|w104|w063|w038|w105|w066|w106|w042;
	wire x029 = w107|w050|w108|w109|w110|w111|w112|w113;
	wire x030 = w114|w115|w116|w117|w118|w119|w120|w121|w122;
	wire x031 = w045|w046|w028|w048|w031;
	wire x032 = w123|w124|w125|w126|w127|w058|w034;
	wire x033 = w128|w075|w129|w130;
	wire x034 = w016|w017|w131|w132|w133|w134|w135|w136|w137|w138|w019|w020|w021|w022|w139|w025|w140;
	wire x035 = w141|w142|w143|w144|w145|w146|w007|w147|w034;
	wire x036 = w148;
	wire x037 = w033;
	wire x038 = w092|w124|w027|w019|w149|w021|w033|w034;
	wire x039 = w092|w027|w019|w149|w021|w033|w034;
	wire x040 = w091|w150|w038|w151|w033|w042;
	wire x041 = w152|w153|w154|w155|w033|w112;
	wire x042 = w156|w027|w016|w157|w158|w159|w007|w020|w032|w160|w161|w162|w163;
	wire x043 = w035|w036|w037|w040|w164|w041|w165|w033|w042;
	wire x044 = w166|w036|w029|w019|w164|w032|w167|w021|w034|w162;
	wire x045 = w168|w169|w043|w074|w048|w049;
	wire x046 = w170|w171|w172|w161|w025;
	wire x047 = w173|w174|w175;
	wire x048 = w176;
	wire x049 = w177;
	wire x050 = w178|w179;
	wire x051 = w180;
	wire x052 = w181|w182;
	wire x053 = w183;
	wire x054 = w184|w062|w185|w070|w146|w186|w187;
	wire x055 = w188|w189|w190|w191|w192|w193|w194|w195|w196;
	wire x056 = w197|w198|w199|w200|w201|w202;
	wire x057 = w043;
	wire x058 = w028|w074;
	wire x059 = w203|w204|w205|w206;
	wire x060 = w207|w208|w209|w210|w211;
	wire x061 = w175|w062|w185|w038|w212|w213;
	wire x062 = w188|w214|w215|w216|w217|w218|w219|w195;
	wire x063 = w198|w220|w126|w221|w201;
	wire x064 = w203|w222|w223|w224|w118|w225;
	wire x065 = w028;
	wire x066 = w209|w226|w227|w228|w229;
	wire x067 = w062|w185|w230|w038|w231|w213;
	wire x068 = w215|w216|w190|w232|w233|w234|w235|w236;
	wire x069 = w198|w220|w237|w238|w239|w240;
	wire x070 = w028|w241;
	wire x071 = w203|w204|w242|w118|w243;
	wire x072 = w209|w244|w245;
	wire x073 = w246|w173|w174;
	wire x074 = w247|w176|w248;
	wire x075 = w178;
	wire x076 = w249|w177|w250;
	wire x077 = w251;
	wire x078 = w252;
	wire x079 = w253|w062|w254|w255;
	wire x080 = w028|w031;
	wire x081 = w198|w193;
	wire x082 = w256|w062|w185|w257|w200|w258|w254;
	wire x083 = w259|w043|w260|w261|w044;
	wire x084 = w262|w263|w028|w264|w265|w266|w267|w031;
	wire x085 = w178|w268|w269|w270;
	wire x086 = w047|w259|w060|w146|w044;
	wire x087 = w271|w272|w273|w274|w185|w275|w276;
	wire x088 = w277|w278|w028|w071|w072|w031;
	wire x089 = w279|w280|w281|w089|w025;
	wire x090 = w068|w282|w283|w284;
	wire x091 = w059|w260;
	wire x092 = w285|w257;
	wire x093 = w286|w287|w288|w289;
	wire x094 = w290|w282|w291|w265|w283;
	wire x095 = w292;
	wire x096 = w287|w288|w070|w030;
	wire x097 = w293|w056|w057;
	wire x098 = w294|w295|w064;
	wire x099 = w208|w076;
	wire x100 = w296;
	wire x101 = w297;
	wire x102 = w144|w152|w146|w298|w155|w014|w034;
	wire x103 = w092|w027|w019|w149|w021|w034;
	wire x104 = w084|w299|w089|w014|w300;
	wire x105 = w301|w302|w303|w304|w305;
	wire x106 = w092|w306|w126|w221|w307|w149|w308;
	wire x107 = w097|w099|w165;
	wire x108 = w309;
	wire x109 = w310|w197;
	wire x110 = w311|w312|w184|w313;
	wire x111 = w314;
	wire x112 = w315|w316|w317|w318;
	wire x113 = w319|w077;
	wire x114 = w320;
	wire x115 = w321|w322;
	wire x116 = w323|w324|w320;
	wire x117 = w286|w314;
	wire x118 = w325|w311|w312;
	wire x119 = w310;
	wire x120 = w326;
	wire x121 = w327;
	wire x122 = w328;
	wire x123 = w329|w050;
	wire x124 = w329;
	wire x125 = w330|w053;
	wire x126 = w331;
	wire x127 = w332;
	wire x128 = w333|w334|w335;
	wire x129 = w336;
	wire x130 = w337|w338;
	wire x131 = w339|w340;
	wire x132 = w341;
	wire x133 = w342;
	wire x134 = w343;
	wire x135 = w344|w333|w334;
	wire x136 = w345|w341|w346;
	wire x137 = w347|w343|w348;
	wire x138 = w337;
	wire x139 = w349;
	wire x140 = w350;
	wire x141 = w351;
	wire x142 = w352;
	wire x143 = w353|w354;
	wire x144 = w355|w356|w357;
	wire x145 = w358;
	wire x146 = w359|w360;
	wire x147 = w361;
	wire x148 = w362;
	wire x149 = w363;
	wire x150 = w364|w355|w356;
	wire x151 = w365|w366|w361;
	wire x152 = w367;
	wire x153 = w368|w362;
	wire x154 = w359;
	wire x155 = w215|w217|w218;
	wire x156 = w226;
	wire x157 = w222|w131;
	wire x158 = w126|w369;
	wire x159 = w038;
	wire x160 = w370;
	wire x161 = w371;
	wire x162 = w317|w318;
	wire x163 = w313;
	wire x164 = w322;
	wire x165 = w372|w373;
	wire x166 = w374|w375|w376;
	wire x167 = w377;
	wire x168 = w378|w379;
	wire x169 = w380|w381|w382;
	wire x170 = w383|w384;
	wire x171 = w385|w386;
	wire x172 = w387;
	wire x173 = w388|w389|w390;
	wire x174 = w391|w392|w393;
	wire x175 = w394|w395;
	wire x176 = w396;
	wire x177 = w397|w376;
	wire x178 = w398|w399;
	wire x179 = w400;
	wire x180 = w242|w205|w401|w402;
	wire x181 = w403;
	wire x182 = w404;
	wire x183 = w405|w406|w401|w395|w407;
	wire x184 = w408|w409;
	wire x185 = w410;
	wire x186 = w411;
	wire x187 = w412;
	wire x188 = w413;
	wire x189 = w414;
	wire x190 = w415;
	wire x191 = w416|w417;
	wire x192 = w387|w418|w419|w420;
	wire x193 = w392|w393|w421;
	wire x194 = w422|w223;
	wire x195 = w390|w423;
	wire x196 = w386;
	wire x197 = w193;
	wire x198 = w199|w200;
	wire x199 = w146;
	wire x200 = w424|w425|w231;
	wire x201 = w426|w238|w239;
	wire x202 = w427|w241;
	wire x203 = w428;
	wire x204 = w234;
	wire x205 = w429;
	wire x206 = w430;
	wire x207 = w234|w431|w432;
	wire x208 = w231|w433;
	wire x209 = w241;
	wire x210 = w238|w239|w434;
	wire x211 = w435;
	wire x212 = w436;
	wire x213 = w437;
	wire x214 = w438;
	
	wire y000 = (t0)|(t1 & x001)|(t2 & x000)|(t3 & x002)|(t4 & x003)|(t5 & x005)|(t6 & x004);
	wire y001 = (t2 & x007)|(t3 & x006)|(t4 & x008)|(t5 & x009);
	wire y002 = (t1 & x016)|(t2 & x015)|(t3 & x010)|(t4 & x012)|(t5 & x013)|(t6 & x011)|(t7 & x014);
	wire y003 = (t2 & x017)|(t3 & x018);
	wire y004 = (t2 & x019)|(t3 & x020)|(t4 & x020);
	wire y005 = (t2 & x017);
	wire y006 = (t3 & x017)|(t4 & x018);
	wire y007 = (t2 & x021)|(t4 & x017);
	wire y008 = (t5 & x017);
	wire y009 = (t1 & x022)|(t3 & x023)|(t5 & x017);
	wire y010 = (t6 & x017);
	wire y011 = (t2 & x024)|(t3 & x025)|(t4 & x023)|(t5 & x018)|(t6 & x017);
	wire y012 = (t2 & x026)|(t4 & x027)|(t5 & x018)|(t6 & x017);
	wire y013 = (t1 & x030)|(t2 & x033)|(t3 & x029)|(t4 & x032)|(t5 & x028)|(t6 & x031)|(t7 & x004);
	wire y014 = (t1 & x034)|(t2 & x035)|(t5 & x036);
	wire y015 = (t1 & x037);
	wire y016 = (t1 & x038)|(t2 & x025);
	wire y017 = (t2 & x037)|(t3 & x023)|(t4 & x023);
	wire y018 = (t2 & x039)|(t3 & x040);
	wire y019 = (t2 & x041);
	wire y020 = (t2 & x037);
	wire y021 = (t3 & x023);
	wire y022 = (t2 & x046)|(t3 & x042)|(t4 & x044)|(t5 & x043)|(t6 & x045)|(t7 & x004);
	wire y023 = (t1 & x051)|(t2 & x053)|(t3 & x052)|(t4 & x050)|(t5 & x047)|(t6 & x048)|(t7 & x049);
	wire y024 = (t1 & x059)|(t2 & x060)|(t3 & x055)|(t4 & x056)|(t5 & x054)|(t6 & x058)|(t7 & x057);
	wire y025 = (t1 & x064)|(t2 & x066)|(t3 & x062)|(t4 & x063)|(t5 & x061)|(t6 & x065)|(t7 & x057);
	wire y026 = (t1 & x071)|(t2 & x072)|(t3 & x068)|(t4 & x069)|(t5 & x067)|(t6 & x070)|(t7 & x057);
	wire y027 = (t1 & x077)|(t2 & x075)|(t3 & x073)|(t4 & x074)|(t5 & x076)|(t6 & x078);
	wire y028 = (t2 & x081)|(t3 & x079)|(t4 & x080)|(t5 & x004);
	wire y029 = (t2 & x081)|(t3 & x082)|(t4 & x084)|(t5 & x083);
	wire y030 = (t3 & x085)|(t4 & x087)|(t5 & x088)|(t6 & x086)|(t7 & x014);
	wire y031 = (t1 & x089);
	wire y032 = (t2 & x092)|(t3 & x090)|(t4 & x091);
	wire y033 = (t3 & x092)|(t4 & x094)|(t5 & x093)|(t6 & x095);
	wire y034 = (t1 & x016)|(t2 & x099)|(t3 & x097)|(t4 & x098)|(t5 & x096)|(t6 & x095);
	wire y035 = (t1 & x100);
	wire y036 = (t1 & x101);
	wire y038 = (t1 & x101)|(t2 & x102)|(t3 & x025);
	wire y041 = (t2 & x101)|(t3 & x103)|(t4 & x025);
	wire y042 = (t2 & x101);
	wire y044 = (t2 & x101)|(t3 & x101);
	wire y046 = (t2 & x104);
	wire y047 = (t2 & x025);
	wire y048 = (t2 & x105)|(t3 & x025);
	wire y049 = (t2 & x106)|(t3 & x107);
	wire y050 = (t1 & x108);
	wire y051 = (t1 & x113)|(t2 & x115)|(t3 & x112)|(t4 & x109)|(t5 & x110)|(t6 & x114)|(t7 & x111);
	wire y052 = (t1 & x120)|(t2 & x119)|(t3 & x118)|(t4 & x116)|(t5 & x117);
	wire y053 = (t2 & x121)|(t3 & x122);
	wire y054 = (t2 & x123)|(t3 & x124)|(t4 & x009);
	wire y055 = (t3 & x125);
	wire y056 = (t1 & x126);
	wire y057 = (t1 & x127);
	wire y058 = (t3 & x036)|(t4 & x009);
	wire y059 = (t4 & x036)|(t5 & x009);
	wire y060 = (t1 & x129)|(t2 & x133)|(t3 & x131)|(t4 & x130)|(t5 & x128)|(t6 & x134)|(t7 & x132);
	wire y061 = (t1 & x139)|(t2 & x138)|(t3 & x135)|(t4 & x137)|(t5 & x136)|(t6 & x140);
	wire y062 = (t1 & x141);
	wire y063 = (t1 & x142);
	wire y064 = (t1 & x149)|(t2 & x145)|(t3 & x143)|(t4 & x146)|(t5 & x144)|(t6 & x147)|(t7 & x148);
	wire y065 = (t1 & x152)|(t2 & x154)|(t3 & x150)|(t4 & x151)|(t5 & x153);
	wire y066 = (t1 & x157)|(t2 & x156)|(t3 & x155)|(t4 & x158)|(t5 & x159);
	wire y067 = (t2 & x027);
	wire y068 = (t1 & x160);
	wire y069 = (t1 & x161);
	wire y070 = (t1 & x016)|(t2 & x164)|(t3 & x162)|(t5 & x163);
	wire y072 = (t1 & x166)|(t2 & x167)|(t3 & x165);
	wire y073 = (t1 & x170)|(t2 & x168)|(t3 & x169);
	wire y074 = (t1 & x175)|(t2 & x172)|(t3 & x174)|(t4 & x173)|(t5 & x171);
	wire y075 = (t1 & x177)|(t2 & x176)|(t3 & x178)|(t4 & x179);
	wire y076 = (t1 & x180);
	wire y077 = (t1 & x181);
	wire y078 = (t1 & x182);
	wire y079 = (t1 & x183)|(t2 & x186)|(t3 & x184)|(t4 & x185)|(t5 & x187);
	wire y080 = (t1 & x188);
	wire y081 = (t1 & x189);
	wire y082 = (t1 & x190);
	wire y083 = (t1 & x194)|(t2 & x191)|(t3 & x192)|(t4 & x193)|(t5 & x195)|(t6 & x196);
	wire y084 = (t3 & x197)|(t4 & x198)|(t5 & x199)|(t6 & x014);
	wire y085 = (t1 & x203)|(t2 & x204)|(t3 & x201)|(t4 & x200)|(t5 & x202);
	wire y086 = (t1 & x205);
	wire y087 = (t1 & x206);
	wire y088 = (t1 & x211)|(t2 & x212)|(t3 & x207)|(t4 & x210)|(t5 & x208)|(t6 & x209);
	wire y089 = (t1 & x213);
	wire y090 = (t1 & x214);
	wire y091 = (t0);
	
	assign O_control[  0] = y000;
	assign O_control[  1] = y001;
	assign O_control[  2] = y002;
	assign O_control[  3] = y003;
	assign O_control[  4] = y004;
	assign O_control[  5] = y005;
	assign O_control[  6] = y006;
	assign O_control[  7] = y007;
	assign O_control[  8] = y008;
	assign O_control[  9] = y009;
	assign O_control[ 10] = y010;
	assign O_control[ 11] = y011;
	assign O_control[ 12] = y012;
	assign O_control[ 13] = y013;
	assign O_control[ 14] = y014;
	assign O_control[ 15] = y015;
	assign O_control[ 16] = y016;
	assign O_control[ 17] = y017;
	assign O_control[ 18] = y018;
	assign O_control[ 19] = y019;
	assign O_control[ 20] = y020;
	assign O_control[ 21] = y021;
	assign O_control[ 22] = y022;
	assign O_control[ 23] = y023;
	assign O_control[ 24] = y024;
	assign O_control[ 25] = y025;
	assign O_control[ 26] = y026;
	assign O_control[ 27] = y027;
	assign O_control[ 28] = y028;
	assign O_control[ 29] = y029;
	assign O_control[ 30] = y030;
	assign O_control[ 31] = y031;
	assign O_control[ 32] = y032;
	assign O_control[ 33] = y033;
	assign O_control[ 34] = y034;
	assign O_control[ 35] = y035;
	assign O_control[ 36] = y036;
	assign O_control[ 37] = y036;
	assign O_control[ 38] = y038;
	assign O_control[ 39] = y036;
	assign O_control[ 40] = y036;
	assign O_control[ 41] = y041;
	assign O_control[ 42] = y042;
	assign O_control[ 43] = y041;
	assign O_control[ 44] = y044;
	assign O_control[ 45] = y042;
	assign O_control[ 46] = y046;
	assign O_control[ 47] = y047;
	assign O_control[ 48] = y048;
	assign O_control[ 49] = y049;
	assign O_control[ 50] = y050;
	assign O_control[ 51] = y051;
	assign O_control[ 52] = y052;
	assign O_control[ 53] = y053;
	assign O_control[ 54] = y054;
	assign O_control[ 55] = y055;
	assign O_control[ 56] = y056;
	assign O_control[ 57] = y057;
	assign O_control[ 58] = y058;
	assign O_control[ 59] = y059;
	assign O_control[ 60] = y060;
	assign O_control[ 61] = y061;
	assign O_control[ 62] = y062;
	assign O_control[ 63] = y063;
	assign O_control[ 64] = y064;
	assign O_control[ 65] = y065;
	assign O_control[ 66] = y066;
	assign O_control[ 67] = y067;
	assign O_control[ 68] = y068;
	assign O_control[ 69] = y069;
	assign O_control[ 70] = y070;
	assign O_control[ 71] = y070;
	assign O_control[ 72] = y072;
	assign O_control[ 73] = y073;
	assign O_control[ 74] = y074;
	assign O_control[ 75] = y075;
	assign O_control[ 76] = y076;
	assign O_control[ 77] = y077;
	assign O_control[ 78] = y078;
	assign O_control[ 79] = y079;
	assign O_control[ 80] = y080;
	assign O_control[ 81] = y081;
	assign O_control[ 82] = y082;
	assign O_control[ 83] = y083;
	assign O_control[ 84] = y084;
	assign O_control[ 85] = y085;
	assign O_control[ 86] = y086;
	assign O_control[ 87] = y087;
	assign O_control[ 88] = y088;
	assign O_control[ 89] = y089;
	assign O_control[ 90] = y090;
	assign O_control[ 91] = y091;
	assign O_control[ 92] = y091;
endmodule