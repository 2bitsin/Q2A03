
module core_decoder(I_ir, I_t, O_control);
	input wire[7:0] I_ir;
	input wire[3:0] I_t;
	output wire[94:0] O_control;
	
	wire w000 = (I_ir ==? 8'b0??11??1);
	wire w001 = (I_ir ==? 8'b0???11??);
	wire w002 = (I_ir ==? 8'b11?11?11);
	wire w003 = (I_ir ==? 8'b1?1?11??);
	wire w004 = (I_ir ==? 8'b1??011??);
	wire w005 = (I_ir ==? 8'b?1??11??);
	wire w006 = (I_ir ==? 8'b???11?01);
	wire w007 = (I_ir ==? 8'b0??1???1);
	wire w008 = (I_ir ==? 8'b0???0??1);
	wire w009 = (I_ir ==? 8'b0????1??);
	wire w010 = (I_ir ==? 8'b11000?1?);
	wire w011 = (I_ir ==? 8'b11??0??1);
	wire w012 = (I_ir ==? 8'b11??1???);
	wire w013 = (I_ir ==? 8'b1?10????);
	wire w014 = (I_ir ==? 8'b1?110??1);
	wire w015 = (I_ir ==? 8'b1?1111??);
	wire w016 = (I_ir ==? 8'b???00??1);
	wire w017 = (I_ir ==? 8'b???0111?);
	wire w018 = (I_ir ==? 8'b???0??0?);
	wire w019 = (I_ir ==? 8'b???11101);
	wire w020 = (I_ir ==? 8'b????01??);
	wire w021 = (I_ir ==? 8'b????10?0);
	wire w022 = (I_ir ==? 8'b?????00?);
	wire w023 = (I_ir ==? 8'b0?100000);
	wire w024 = (I_ir ==? 8'b0?101?00);
	wire w025 = (I_ir ==? 8'b0??0000?);
	wire w026 = (I_ir ==? 8'b0???0?11);
	wire w027 = (I_ir ==? 8'b0????110);
	wire w028 = (I_ir ==? 8'b1001??01);
	wire w029 = (I_ir ==? 8'b11?011??);
	wire w030 = (I_ir ==? 8'b?0?000?1);
	wire w031 = (I_ir ==? 8'b?0?011??);
	wire w032 = (I_ir ==? 8'b?0??0001);
	wire w033 = (I_ir ==? 8'b?1?011?1);
	wire w034 = (I_ir ==? 8'b?1?0?11?);
	wire w035 = (I_ir ==? 8'b?1??00?1);
	wire w036 = (I_ir ==? 8'b?1???110);
	wire w037 = (I_ir ==? 8'b??1?00?1);
	wire w038 = (I_ir ==? 8'b???101??);
	wire w039 = (I_ir ==? 8'b0??0??00);
	wire w040 = (I_ir ==? 8'b101?0??1);
	wire w041 = (I_ir ==? 8'b?1?111??);
	wire w042 = (I_ir ==? 8'b?1?1???1);
	wire w043 = (I_ir ==? 8'b??1111??);
	wire w044 = (I_ir ==? 8'b???0?1??);
	wire w045 = (I_ir ==? 8'b???1??01);
	wire w046 = (I_ir ==? 8'b011?11?0);
	wire w047 = (I_ir ==? 8'b0??111??);
	wire w048 = (I_ir ==? 8'b0??11?11);
	wire w049 = (I_ir ==? 8'b0????11?);
	wire w050 = (I_ir ==? 8'b100?0001);
	wire w051 = (I_ir ==? 8'b?1?11?11);
	wire w052 = (I_ir ==? 8'b?1???11?);
	wire w053 = (I_ir ==? 8'b???000?1);
	wire w054 = (I_ir ==? 8'b0??1?11?);
	wire w055 = (I_ir ==? 8'b0??1??11);
	wire w056 = (I_ir ==? 8'b0???111?);
	wire w057 = (I_ir ==? 8'b101?00?1);
	wire w058 = (I_ir ==? 8'b11?1?011);
	wire w059 = (I_ir ==? 8'b?1?1?11?);
	wire w060 = (I_ir ==? 8'b?1??111?);
	wire w061 = (I_ir ==? 8'b????0001);
	wire w062 = (I_ir ==? 8'b0???0011);
	wire w063 = (I_ir ==? 8'b?1??0011);
	wire w064 = (I_ir ==? 8'b00000000);
	wire w065 = (I_ir ==? 8'b00?1111?);
	wire w066 = (I_ir ==? 8'b00??0011);
	wire w067 = (I_ir ==? 8'b?1?1111?);
	wire w068 = (I_ir ==? 8'b?1?1?011);
	wire w069 = (I_ir ==? 8'b0?101000);
	wire w070 = (I_ir ==? 8'b0??00000);
	wire w071 = (I_ir ==? 8'b0??0?000);
	wire w072 = (I_ir ==? 8'b01000000);
	wire w073 = (I_ir ==? 8'b00?00000);
	wire w074 = (I_ir ==? 8'b0??0011?);
	wire w075 = (I_ir ==? 8'b100011??);
	wire w076 = (I_ir ==? 8'b100101??);
	wire w077 = (I_ir ==? 8'b?1?0011?);
	wire w078 = (I_ir ==? 8'b0??11110);
	wire w079 = (I_ir ==? 8'b11?1111?);
	wire w080 = (I_ir ==? 8'b00?0?110);
	wire w081 = (I_ir ==? 8'b0??01111);
	wire w082 = (I_ir ==? 8'b0??1011?);
	wire w083 = (I_ir ==? 8'b10011?01);
	wire w084 = (I_ir ==? 8'b11??011?);
	wire w085 = (I_ir ==? 8'b?1?0111?);
	wire w086 = (I_ir ==? 8'b?1??0110);
	wire w087 = (I_ir ==? 8'b00?10110);
	wire w088 = (I_ir ==? 8'b0???1110);
	wire w089 = (I_ir ==? 8'b100000?1);
	wire w090 = (I_ir ==? 8'b11?1?11?);
	wire w091 = (I_ir ==? 8'b11??111?);
	wire w092 = (I_ir ==? 8'b?1?1?110);
	wire w093 = (I_ir ==? 8'b11??0011);
	wire w094 = (I_ir ==? 8'b0?001000);
	wire w095 = (I_ir ==? 8'b100001??);
	wire w096 = (I_ir ==? 8'b11001011);
	wire w097 = (I_ir ==? 8'b00100000);
	wire w098 = (I_ir ==? 8'b0000?000);
	wire w099 = (I_ir ==? 8'b00001000);
	wire w100 = (I_ir ==? 8'b00100?00);
	wire w101 = (I_ir ==? 8'b001011??);
	wire w102 = (I_ir ==? 8'b0?00?1??);
	wire w103 = (I_ir ==? 8'b0??10??1);
	wire w104 = (I_ir ==? 8'b11010??1);
	wire w105 = (I_ir ==? 8'b?0?10001);
	wire w106 = (I_ir ==? 8'b?110?11?);
	wire w107 = (I_ir ==? 8'b??110??1);
	wire w108 = (I_ir ==? 8'b???0?1?1);
	wire w109 = (I_ir ==? 8'b01101100);
	wire w110 = (I_ir ==? 8'b00?11??1);
	wire w111 = (I_ir ==? 8'b0?0?11??);
	wire w112 = (I_ir ==? 8'b0?1?11?1);
	wire w113 = (I_ir ==? 8'b?01?11??);
	wire w114 = (I_ir ==? 8'b??1?111?);
	wire w115 = (I_ir ==? 8'b0??100?1);
	wire w116 = (I_ir ==? 8'b101100?1);
	wire w117 = (I_ir ==? 8'b?1?100?1);
	wire w118 = (I_ir ==? 8'b???10001);
	wire w119 = (I_ir ==? 8'b01001100);
	wire w120 = (I_ir ==? 8'b0010000?);
	wire w121 = (I_ir ==? 8'b01?0000?);
	wire w122 = (I_ir ==? 8'b0??0111?);
	wire w123 = (I_ir ==? 8'b10?000?1);
	wire w124 = (I_ir ==? 8'b?1?1011?);
	wire w125 = (I_ir ==? 8'b00?0110?);
	wire w126 = (I_ir ==? 8'b10?011??);
	wire w127 = (I_ir ==? 8'b10?101??);
	wire w128 = (I_ir ==? 8'b1??0110?);
	wire w129 = (I_ir ==? 8'b???01101);
	wire w130 = (I_ir ==? 8'b???1010?);
	wire w131 = (I_ir ==? 8'b???10?00);
	wire w132 = (I_ir ==? 8'b1010?0?0);
	wire w133 = (I_ir ==? 8'b10?0?000);
	wire w134 = (I_ir ==? 8'b11?010??);
	wire w135 = (I_ir ==? 8'b11?0?0?0);
	wire w136 = (I_ir ==? 8'b1?1010?1);
	wire w137 = (I_ir ==? 8'b1???10?0);
	wire w138 = (I_ir ==? 8'b???01001);
	wire w139 = (I_ir ==? 8'b???110?0);
	wire w140 = (I_ir ==? 8'b????1010);
	wire w141 = (I_ir ==? 8'b00?0011?);
	wire w142 = (I_ir ==? 8'b011?1100);
	wire w143 = (I_ir ==? 8'b0??1110?);
	wire w144 = (I_ir ==? 8'b101111??);
	wire w145 = (I_ir ==? 8'b11?1110?);
	wire w146 = (I_ir ==? 8'b0100?100);
	wire w147 = (I_ir ==? 8'b10?001??);
	wire w148 = (I_ir ==? 8'b???0010?);
	wire w149 = (I_ir ==? 8'b101010?1);
	wire w150 = (I_ir ==? 8'b11?0?0?1);
	wire w151 = (I_ir ==? 8'b1?10001?);
	wire w152 = (I_ir ==? 8'b1??0000?);
	wire w153 = (I_ir ==? 8'b1??0?1??);
	wire w154 = (I_ir ==? 8'b?01?000?);
	wire w155 = (I_ir ==? 8'b???1000?);
	wire w156 = (I_ir ==? 8'b??????01);
	wire w157 = (I_ir ==? 8'b01??11?1);
	wire w158 = (I_ir ==? 8'b0?0111??);
	wire w159 = (I_ir ==? 8'b0?0?111?);
	wire w160 = (I_ir ==? 8'b110?11??);
	wire w161 = (I_ir ==? 8'b??1?11??);
	wire w162 = (I_ir ==? 8'b01100000);
	wire w163 = (I_ir ==? 8'b?1?11??1);
	wire w164 = (I_ir ==? 8'b0???00?1);
	wire w165 = (I_ir ==? 8'b11??00?1);
	wire w166 = (I_ir ==? 8'b0??1?1??);
	wire w167 = (I_ir ==? 8'b1?11110?);
	wire w168 = (I_ir ==? 8'b1??1?101);
	wire w169 = (I_ir ==? 8'b?1?1?1??);
	wire w170 = (I_ir ==? 8'b00???11?);
	wire w171 = (I_ir ==? 8'b11??11??);
	wire w172 = (I_ir ==? 8'b1?110?11);
	wire w173 = (I_ir ==? 8'b1??1011?);
	wire w174 = (I_ir ==? 8'b??11?1??);
	wire w175 = (I_ir ==? 8'b???10?0?);
	wire w176 = (I_ir ==? 8'b???1?001);
	wire w177 = (I_ir ==? 8'b????1101);
	wire w178 = (I_ir ==? 8'b?1?1??11);
	wire w179 = (I_ir ==? 8'b??1100?1);
	wire w180 = (I_ir ==? 8'b000111??);
	wire w181 = (I_ir ==? 8'b??110011);
	wire w182 = (I_ir ==? 8'b00?11011);
	wire w183 = (I_ir ==? 8'b0??1111?);
	wire w184 = (I_ir ==? 8'b0?010?11);
	wire w185 = (I_ir ==? 8'b?0110?11);
	wire w186 = (I_ir ==? 8'b?1?10?11);
	wire w187 = (I_ir ==? 8'b00001111);
	wire w188 = (I_ir ==? 8'b00010111);
	wire w189 = (I_ir ==? 8'b000?0001);
	wire w190 = (I_ir ==? 8'b00011?11);
	wire w191 = (I_ir ==? 8'b000?0011);
	wire w192 = (I_ir ==? 8'b00000111);
	wire w193 = (I_ir ==? 8'b00011?01);
	wire w194 = (I_ir ==? 8'b00001001);
	wire w195 = (I_ir ==? 8'b00001101);
	wire w196 = (I_ir ==? 8'b00010101);
	wire w197 = (I_ir ==? 8'b00000101);
	wire w198 = (I_ir ==? 8'b001?0001);
	wire w199 = (I_ir ==? 8'b0??10111);
	wire w200 = (I_ir ==? 8'b?11?0001);
	wire w201 = (I_ir ==? 8'b??0?0001);
	wire w202 = (I_ir ==? 8'b0010110?);
	wire w203 = (I_ir ==? 8'b00?01101);
	wire w204 = (I_ir ==? 8'b0??10101);
	wire w205 = (I_ir ==? 8'b100011?1);
	wire w206 = (I_ir ==? 8'b100101?1);
	wire w207 = (I_ir ==? 8'b11?00111);
	wire w208 = (I_ir ==? 8'b?1?01101);
	wire w209 = (I_ir ==? 8'b?1?10101);
	wire w210 = (I_ir ==? 8'b??010101);
	wire w211 = (I_ir ==? 8'b00111?01);
	wire w212 = (I_ir ==? 8'b0??00111);
	wire w213 = (I_ir ==? 8'b11?01111);
	wire w214 = (I_ir ==? 8'b11?10111);
	wire w215 = (I_ir ==? 8'b?1?11?01);
	wire w216 = (I_ir ==? 8'b??011?01);
	wire w217 = (I_ir ==? 8'b0??01001);
	wire w218 = (I_ir ==? 8'b0??01010);
	wire w219 = (I_ir ==? 8'b101010?0);
	wire w220 = (I_ir ==? 8'b11?010?1);
	wire w221 = (I_ir ==? 8'b0010010?);
	wire w222 = (I_ir ==? 8'b01001000);
	wire w223 = (I_ir ==? 8'b0??00101);
	wire w224 = (I_ir ==? 8'b100001?1);
	wire w225 = (I_ir ==? 8'b11?00101);
	wire w226 = (I_ir ==? 8'b?1??0001);
	wire w227 = (I_ir ==? 8'b??1?0001);
	wire w228 = (I_ir ==? 8'b00?10101);
	wire w229 = (I_ir ==? 8'b01101000);
	wire w230 = (I_ir ==? 8'b0??01101);
	wire w231 = (I_ir ==? 8'b101011??);
	wire w232 = (I_ir ==? 8'b101101??);
	wire w233 = (I_ir ==? 8'b11?0110?);
	wire w234 = (I_ir ==? 8'b0??11?01);
	wire w235 = (I_ir ==? 8'b1?111?01);
	wire w236 = (I_ir ==? 8'b101000?0);
	wire w237 = (I_ir ==? 8'b11?00000);
	wire w238 = (I_ir ==? 8'b1?100000);
	wire w239 = (I_ir ==? 8'b?1?01001);
	wire w240 = (I_ir ==? 8'b101001??);
	wire w241 = (I_ir ==? 8'b11?0010?);
	wire w242 = (I_ir ==? 8'b?010010?);
	wire w243 = (I_ir ==? 8'b?1?00101);
	wire w244 = (I_ir ==? 8'b0???0001);
	wire w245 = (I_ir ==? 8'b11111?11);
	wire w246 = (I_ir ==? 8'b101011?1);
	wire w247 = (I_ir ==? 8'b101101?1);
	wire w248 = (I_ir ==? 8'b11100111);
	wire w249 = (I_ir ==? 8'b1?101101);
	wire w250 = (I_ir ==? 8'b??110101);
	wire w251 = (I_ir ==? 8'b101111?1);
	wire w252 = (I_ir ==? 8'b11101111);
	wire w253 = (I_ir ==? 8'b11110111);
	wire w254 = (I_ir ==? 8'b??111?01);
	wire w255 = (I_ir ==? 8'b111?0011);
	wire w256 = (I_ir ==? 8'b10011000);
	wire w257 = (I_ir ==? 8'b?0001010);
	wire w258 = (I_ir ==? 8'b101001?1);
	wire w259 = (I_ir ==? 8'b1?100101);
	wire w260 = (I_ir ==? 8'b00000110);
	wire w261 = (I_ir ==? 8'b0000?110);
	wire w262 = (I_ir ==? 8'b000?0110);
	wire w263 = (I_ir ==? 8'b0001?110);
	wire w264 = (I_ir ==? 8'b000?1110);
	wire w265 = (I_ir ==? 8'b00001010);
	wire w266 = (I_ir ==? 8'b00011110);
	wire w267 = (I_ir ==? 8'b00?10111);
	wire w268 = (I_ir ==? 8'b?1?01111);
	wire w269 = (I_ir ==? 8'b?1?10111);
	wire w270 = (I_ir ==? 8'b0?100110);
	wire w271 = (I_ir ==? 8'b11?00110);
	wire w272 = (I_ir ==? 8'b?1100110);
	wire w273 = (I_ir ==? 8'b0?111110);
	wire w274 = (I_ir ==? 8'b11?11110);
	wire w275 = (I_ir ==? 8'b?1111110);
	wire w276 = (I_ir ==? 8'b0?101110);
	wire w277 = (I_ir ==? 8'b0?110110);
	wire w278 = (I_ir ==? 8'b11?01110);
	wire w279 = (I_ir ==? 8'b11?10110);
	wire w280 = (I_ir ==? 8'b?1101110);
	wire w281 = (I_ir ==? 8'b?1110110);
	wire w282 = (I_ir ==? 8'b0?10011?);
	wire w283 = (I_ir ==? 8'b11?0011?);
	wire w284 = (I_ir ==? 8'b?1?00111);
	wire w285 = (I_ir ==? 8'b0?001111);
	wire w286 = (I_ir ==? 8'b0?10111?);
	wire w287 = (I_ir ==? 8'b0?11011?);
	wire w288 = (I_ir ==? 8'b0?1?0110);
	wire w289 = (I_ir ==? 8'b11?0?11?);
	wire w290 = (I_ir ==? 8'b11?1011?);
	wire w291 = (I_ir ==? 8'b0?11?110);
	wire w292 = (I_ir ==? 8'b0?1?1110);
	wire w293 = (I_ir ==? 8'b00?10??1);
	wire w294 = (I_ir ==? 8'b1??10001);
	wire w295 = (I_ir ==? 8'b?1010??1);
	wire w296 = (I_ir ==? 8'b0??01110);
	wire w297 = (I_ir ==? 8'b?1?01110);
	wire w298 = (I_ir ==? 8'b?1?10110);
	wire w299 = (I_ir ==? 8'b0??00110);
	wire w300 = (I_ir ==? 8'b00111110);
	wire w301 = (I_ir ==? 8'b0?01?110);
	wire w302 = (I_ir ==? 8'b0?0?1110);
	wire w303 = (I_ir ==? 8'b?1?11110);
	wire w304 = (I_ir ==? 8'b0?00?110);
	wire w305 = (I_ir ==? 8'b0??10110);
	wire w306 = (I_ir ==? 8'b0?011110);
	wire w307 = (I_ir ==? 8'b0?000110);
	wire w308 = (I_ir ==? 8'b0?001110);
	wire w309 = (I_ir ==? 8'b0?0?0110);
	wire w310 = (I_ir ==? 8'b00?011??);
	wire w311 = (I_ir ==? 8'b00010000);
	wire w312 = (I_ir ==? 8'b???10000);
	wire w313 = (I_ir ==? 8'b1?11?1??);
	wire w314 = (I_ir ==? 8'b11?10??1);
	wire w315 = (I_ir ==? 8'b???10?01);
	wire w316 = (I_ir ==? 8'b0??110?1);
	wire w317 = (I_ir ==? 8'b1011?11?);
	wire w318 = (I_ir ==? 8'b10?1011?);
	wire w319 = (I_ir ==? 8'b?1?110?1);
	wire w320 = (I_ir ==? 8'b???11001);
	wire w321 = (I_ir ==? 8'b0?01110?);
	wire w322 = (I_ir ==? 8'b?101110?);
	wire w323 = (I_ir ==? 8'b??11110?);
	wire w324 = (I_ir ==? 8'b00011000);
	wire w325 = (I_ir ==? 8'b00100111);
	wire w326 = (I_ir ==? 8'b00101111);
	wire w327 = (I_ir ==? 8'b00110111);
	wire w328 = (I_ir ==? 8'b10000011);
	wire w329 = (I_ir ==? 8'b001?0011);
	wire w330 = (I_ir ==? 8'b00101101);
	wire w331 = (I_ir ==? 8'b00110101);
	wire w332 = (I_ir ==? 8'b10001111);
	wire w333 = (I_ir ==? 8'b10010111);
	wire w334 = (I_ir ==? 8'b00101001);
	wire w335 = (I_ir ==? 8'b00111?11);
	wire w336 = (I_ir ==? 8'b00100101);
	wire w337 = (I_ir ==? 8'b10000111);
	wire w338 = (I_ir ==? 8'b00101110);
	wire w339 = (I_ir ==? 8'b00110110);
	wire w340 = (I_ir ==? 8'b00100110);
	wire w341 = (I_ir ==? 8'b00101010);
	wire w342 = (I_ir ==? 8'b00100100);
	wire w343 = (I_ir ==? 8'b00101100);
	wire w344 = (I_ir ==? 8'b01?00000);
	wire w345 = (I_ir ==? 8'b00101000);
	wire w346 = (I_ir ==? 8'b00110000);
	wire w347 = (I_ir ==? 8'b00111000);
	wire w348 = (I_ir ==? 8'b01001111);
	wire w349 = (I_ir ==? 8'b01010111);
	wire w350 = (I_ir ==? 8'b010?0001);
	wire w351 = (I_ir ==? 8'b01001001);
	wire w352 = (I_ir ==? 8'b01000111);
	wire w353 = (I_ir ==? 8'b01011?01);
	wire w354 = (I_ir ==? 8'b01001101);
	wire w355 = (I_ir ==? 8'b01010101);
	wire w356 = (I_ir ==? 8'b010?0011);
	wire w357 = (I_ir ==? 8'b01000101);
	wire w358 = (I_ir ==? 8'b01011?11);
	wire w359 = (I_ir ==? 8'b01000110);
	wire w360 = (I_ir ==? 8'b0101?110);
	wire w361 = (I_ir ==? 8'b010?1110);
	wire w362 = (I_ir ==? 8'b0100?110);
	wire w363 = (I_ir ==? 8'b010?0110);
	wire w364 = (I_ir ==? 8'b01001010);
	wire w365 = (I_ir ==? 8'b01011110);
	wire w366 = (I_ir ==? 8'b01010000);
	wire w367 = (I_ir ==? 8'b01011000);
	wire w368 = (I_ir ==? 8'b01101101);
	wire w369 = (I_ir ==? 8'b01110101);
	wire w370 = (I_ir ==? 8'b01101111);
	wire w371 = (I_ir ==? 8'b01110111);
	wire w372 = (I_ir ==? 8'b011?0001);
	wire w373 = (I_ir ==? 8'b01100101);
	wire w374 = (I_ir ==? 8'b01100111);
	wire w375 = (I_ir ==? 8'b01111?01);
	wire w376 = (I_ir ==? 8'b01111?11);
	wire w377 = (I_ir ==? 8'b011?0011);
	wire w378 = (I_ir ==? 8'b01101001);
	wire w379 = (I_ir ==? 8'b01100110);
	wire w380 = (I_ir ==? 8'b01101110);
	wire w381 = (I_ir ==? 8'b01110110);
	wire w382 = (I_ir ==? 8'b01101010);
	wire w383 = (I_ir ==? 8'b01111110);
	wire w384 = (I_ir ==? 8'b10111?01);
	wire w385 = (I_ir ==? 8'b01110000);
	wire w386 = (I_ir ==? 8'b01111000);
	wire w387 = (I_ir ==? 8'b10010100);
	wire w388 = (I_ir ==? 8'b1?001100);
	wire w389 = (I_ir ==? 8'b100?1000);
	wire w390 = (I_ir ==? 8'b1100?000);
	wire w391 = (I_ir ==? 8'b1?001000);
	wire w392 = (I_ir ==? 8'b1?000100);
	wire w393 = (I_ir ==? 8'b10000110);
	wire w394 = (I_ir ==? 8'b11100100);
	wire w395 = (I_ir ==? 8'b10001110);
	wire w396 = (I_ir ==? 8'b10010110);
	wire w397 = (I_ir ==? 8'b11101100);
	wire w398 = (I_ir ==? 8'b1110?000);
	wire w399 = (I_ir ==? 8'b1?001010);
	wire w400 = (I_ir ==? 8'b11011110);
	wire w401 = (I_ir ==? 8'b110?0011);
	wire w402 = (I_ir ==? 8'b11000111);
	wire w403 = (I_ir ==? 8'b11001110);
	wire w404 = (I_ir ==? 8'b11010110);
	wire w405 = (I_ir ==? 8'b11011?11);
	wire w406 = (I_ir ==? 8'b11000110);
	wire w407 = (I_ir ==? 8'b11001111);
	wire w408 = (I_ir ==? 8'b11010111);
	wire w409 = (I_ir ==? 8'b10001000);
	wire w410 = (I_ir ==? 8'b11001010);
	wire w411 = (I_ir ==? 8'b10100100);
	wire w412 = (I_ir ==? 8'b1010?000);
	wire w413 = (I_ir ==? 8'b10101100);
	wire w414 = (I_ir ==? 8'b10110100);
	wire w415 = (I_ir ==? 8'b10111100);
	wire w416 = (I_ir ==? 8'b101?1010);
	wire w417 = (I_ir ==? 8'b10?01010);
	wire w418 = (I_ir ==? 8'b10010000);
	wire w419 = (I_ir ==? 8'b10011010);
	wire w420 = (I_ir ==? 8'b1010101?);
	wire w421 = (I_ir ==? 8'b1010?010);
	wire w422 = (I_ir ==? 8'b11101000);
	wire w423 = (I_ir ==? 8'b1010111?);
	wire w424 = (I_ir ==? 8'b1011011?);
	wire w425 = (I_ir ==? 8'b1011111?);
	wire w426 = (I_ir ==? 8'b1010011?);
	wire w427 = (I_ir ==? 8'b101?0011);
	wire w428 = (I_ir ==? 8'b10110000);
	wire w429 = (I_ir ==? 8'b10111000);
	wire w430 = (I_ir ==? 8'b10111010);
	wire w431 = (I_ir ==? 8'b1100010?);
	wire w432 = (I_ir ==? 8'b11?00100);
	wire w433 = (I_ir ==? 8'b1100110?);
	wire w434 = (I_ir ==? 8'b11010101);
	wire w435 = (I_ir ==? 8'b11?01100);
	wire w436 = (I_ir ==? 8'b11011?01);
	wire w437 = (I_ir ==? 8'b11001001);
	wire w438 = (I_ir ==? 8'b110?0001);
	wire w439 = (I_ir ==? 8'b11101110);
	wire w440 = (I_ir ==? 8'b11110110);
	wire w441 = (I_ir ==? 8'b11100110);
	wire w442 = (I_ir ==? 8'b11111110);
	wire w443 = (I_ir ==? 8'b11?01000);
	wire w444 = (I_ir ==? 8'b11010000);
	wire w445 = (I_ir ==? 8'b11011000);
	wire w446 = (I_ir ==? 8'b11101101);
	wire w447 = (I_ir ==? 8'b11110101);
	wire w448 = (I_ir ==? 8'b111?0001);
	wire w449 = (I_ir ==? 8'b11111?01);
	wire w450 = (I_ir ==? 8'b111010?1);
	wire w451 = (I_ir ==? 8'b11100101);
	wire w452 = (I_ir ==? 8'b11110000);
	wire w453 = (I_ir ==? 8'b11111000);
	
	assign O_control[  0] = (((I_t == 4'd2)&(w000|w001|w002|w003|w004|w005|w006))
	                        |((I_t == 4'd1)&(w007|w008|w009|w010|w011|w012|w013|w014|w015|w016|w017|w018|w019|w020|w021|w022))
	                        |((I_t == 4'd5)&(w023))
	                        |((I_t == 4'd0)));
	
	assign O_control[  1] = (((I_t == 4'd2)&(w024|w025|w026|w027|w028|w029|w030|w031|w032|w033|w034|w035|w036|w037|w038))
	                        |((I_t == 4'd1)&(w039|w007|w009|w040|w041|w042|w043|w016|w044|w045|w020))
	                        |((I_t == 4'd3)&(w046|w025|w047|w048|w049|w050|w041|w051|w052|w043|w053|w006))
	                        |((I_t == 4'd4)&(w025|w054|w055|w056|w057|w058|w059|w060|w053|w061))
	                        |((I_t == 4'd6)&(w062|w063))
	                        |((I_t == 4'd5)&(w064|w065|w066|w048|w067|w068|w063))
	                        |((I_t == 4'd0)));
	
	assign O_control[  2] = (((I_t == 4'd3)&(w069|w070))
	                        |((I_t == 4'd2)&(w071))
	                        |((I_t == 4'd4)&(w070))
	                        |((I_t == 4'd5)&(w072)));
	
	assign O_control[  3] = (((I_t == 4'd3)&(w073|w074|w075|w076|w077))
	                        |((I_t == 4'd6)&(w066|w078|w079|w058|w063))
	                        |((I_t == 4'd4)&(w073|w080|w081|w082|w083|w084|w085|w086))
	                        |((I_t == 4'd5)&(w087|w048|w088|w089|w050|w090|w091|w051|w092))
	                        |((I_t == 4'd7)&(w093))
	                        |((I_t == 4'd2)&(w064|w094|w095))
	                        |((I_t == 4'd1)&(w096)));
	
	assign O_control[  4] = (((I_t == 4'd2)&(w064))
	                        |((I_t == 4'd3)&(w097)));
	
	assign O_control[  5] = (((I_t == 4'd2)&(w098|w094))
	                        |((I_t == 4'd3)&(w073))
	                        |((I_t == 4'd4)&(w073)));
	
	assign O_control[  6] = (((I_t == 4'd2)&(w064)));
	
	assign O_control[  7] = (((I_t == 4'd3)&(w064))
	                        |((I_t == 4'd4)&(w097)));
	
	assign O_control[  8] = (((I_t == 4'd2)&(w099))
	                        |((I_t == 4'd4)&(w064)));
	
	assign O_control[  9] = (((I_t == 4'd5)&(w064)));
	
	assign O_control[ 10] = (((I_t == 4'd1)&(w100|w101|w102|w103|w104|w004|w105|w106|w107|w108|w020))
	                        |((I_t == 4'd3)&(w109|w053))
	                        |((I_t == 4'd5)&(w064)));
	
	assign O_control[ 11] = (((I_t == 4'd6)&(w064)));
	
	assign O_control[ 12] = (((I_t == 4'd2)&(w110|w111|w112|w004|w113|w041|w051|w114|w006))
	                        |((I_t == 4'd3)&(w115|w116|w117|w118))
	                        |((I_t == 4'd4)&(w109|w053))
	                        |((I_t == 4'd6)&(w064))
	                        |((I_t == 4'd5)&(w097)));
	
	assign O_control[ 13] = (((I_t == 4'd5)&(w097))
	                        |((I_t == 4'd6)&(w064))
	                        |((I_t == 4'd2)&(w119))
	                        |((I_t == 4'd4)&(w109)));
	
	assign O_control[ 14] = (((I_t == 4'd5)&(w120|w121|w122|w082|w057|w123|w085|w124|w061))
	                        |((I_t == 4'd3)&(w125|w069|w126|w127|w128|w129|w130|w131))
	                        |((I_t == 4'd1)&(w132|w133|w134|w135|w136|w137|w138|w139|w140))
	                        |((I_t == 4'd6)&(w064|w065|w048|w067|w051))
	                        |((I_t == 4'd4)&(w141|w142|w143|w144|w145|w077|w006))
	                        |((I_t == 4'd7)&(w062|w063))
	                        |((I_t == 4'd2)&(w146|w094|w147|w148)));
	
	assign O_control[ 15] = (((I_t == 4'd1)&(w007|w009|w149|w010|w150|w151|w014|w152|w153|w154|w041|w042|w043|w016|w155|w020|w156))
	                        |((I_t == 4'd2)&(w157|w158|w159|w000|w160|w002|w031|w161|w006))
	                        |((I_t == 4'd5)&(w162)));
	
	assign O_control[ 16] = (((I_t == 4'd1)&(w053)));
	
	assign O_control[ 17] = (((I_t == 4'd1)&(w110|w142|w047|w041|w163|w043|w053|w006))
	                        |((I_t == 4'd2)&(w115|w116|w117|w118)));
	
	assign O_control[ 18] = (((I_t == 4'd2)&(w053))
	                        |((I_t == 4'd3)&(w109|w053))
	                        |((I_t == 4'd4)&(w109|w053)));
	
	assign O_control[ 19] = (((I_t == 4'd2)&(w110|w047|w041|w163|w043|w053|w006))
	                        |((I_t == 4'd3)&(w109|w164|w057|w165|w053|w061)));
	
	assign O_control[ 20] = (((I_t == 4'd2)&(w166|w167|w168|w169|w053|w130)));
	
	assign O_control[ 21] = (((I_t == 4'd2)&(w053)));
	
	assign O_control[ 22] = (((I_t == 4'd3)&(w109|w053)));
	
	assign O_control[ 23] = (((I_t == 4'd3)&(w170|w047|w007|w171|w172|w173|w031|w042|w052|w174|w175|w176|w177))
	                        |((I_t == 4'd5)&(w054|w055|w056|w059|w178|w060|w179|w053|w061))
	                        |((I_t == 4'd4)&(w180|w055|w049|w041|w178|w052|w181|w043|w006|w176))
	                        |((I_t == 4'd6)&(w182|w183|w062|w093|w067|w068))
	                        |((I_t == 4'd2)&(w184|w185|w186|w175|w020))
	                        |((I_t == 4'd7)&(w062|w063)));
	
	assign O_control[ 24] = (((I_t == 4'd5)&(w187|w188|w189))
	                        |((I_t == 4'd6)&(w190))
	                        |((I_t == 4'd7)&(w191))
	                        |((I_t == 4'd4)&(w192|w193))
	                        |((I_t == 4'd1)&(w194))
	                        |((I_t == 4'd3)&(w195|w196))
	                        |((I_t == 4'd2)&(w197)));
	
	assign O_control[ 25] = (((I_t == 4'd5)&(w198|w081|w199|w089|w002|w200|w201))
	                        |((I_t == 4'd3)&(w202|w203|w204|w205|w206|w207|w208|w209|w210))
	                        |((I_t == 4'd4)&(w211|w212|w213|w214|w215|w216))
	                        |((I_t == 4'd7)&(w062))
	                        |((I_t == 4'd6)&(w048|w093))
	                        |((I_t == 4'd1)&(w217|w218|w219|w220))
	                        |((I_t == 4'd2)&(w221|w222|w223|w224|w225)));
	
	assign O_control[ 26] = (((I_t == 4'd5)&(w189|w081|w199|w057|w226|w227))
	                        |((I_t == 4'd3)&(w202|w228|w229|w230|w231|w232|w233|w209))
	                        |((I_t == 4'd4)&(w212|w234|w144|w235|w215))
	                        |((I_t == 4'd7)&(w062))
	                        |((I_t == 4'd1)&(w217|w236|w237|w238|w136|w239))
	                        |((I_t == 4'd6)&(w048))
	                        |((I_t == 4'd2)&(w223|w240|w241|w242|w243)));
	
	assign O_control[ 27] = (((I_t == 4'd5)&(w081|w199|w244|w057|w245|w227))
	                        |((I_t == 4'd3)&(w229|w230|w204|w246|w247|w248|w249|w250))
	                        |((I_t == 4'd4)&(w212|w234|w251|w252|w253|w254))
	                        |((I_t == 4'd7)&(w062))
	                        |((I_t == 4'd6)&(w048|w255))
	                        |((I_t == 4'd1)&(w217|w218|w256|w136|w257))
	                        |((I_t == 4'd2)&(w223|w258|w259)));
	
	assign O_control[ 28] = (((I_t == 4'd3)&(w260|w187|w188))
	                        |((I_t == 4'd4)&(w261|w190|w262))
	                        |((I_t == 4'd2)&(w192))
	                        |((I_t == 4'd5)&(w263|w191|w264))
	                        |((I_t == 4'd1)&(w265))
	                        |((I_t == 4'd6)&(w266)));
	
	assign O_control[ 29] = (((I_t == 4'd3)&(w267|w081|w268|w269))
	                        |((I_t == 4'd5)&(w062|w063))
	                        |((I_t == 4'd4)&(w048|w051))
	                        |((I_t == 4'd2)&(w212|w207)));
	
	assign O_control[ 30] = (((I_t == 4'd3)&(w270|w081|w199|w271|w214|w272|w268))
	                        |((I_t == 4'd5)&(w273|w062|w274|w275|w063))
	                        |((I_t == 4'd4)&(w276|w277|w048|w278|w279|w280|w281|w051))
	                        |((I_t == 4'd2)&(w212|w207)));
	
	assign O_control[ 31] = (((I_t == 4'd3)&(w192|w282|w283|w284))
	                        |((I_t == 4'd6)&(w066|w273|w079|w002|w063))
	                        |((I_t == 4'd4)&(w285|w286|w287|w288|w199|w289|w290))
	                        |((I_t == 4'd5)&(w291|w292|w048|w090|w091|w051))
	                        |((I_t == 4'd7)&(w093)));
	
	assign O_control[ 32] = (((I_t == 4'd1)&(w293|w294|w295|w107|w020)));
	
	assign O_control[ 33] = (((I_t == 4'd3)&(w087|w296|w297|w298))
	                        |((I_t == 4'd4)&(w078|w274))
	                        |((I_t == 4'd2)&(w299|w271)));
	
	assign O_control[ 34] = (((I_t == 4'd5)&(w300|w301|w302|w303))
	                        |((I_t == 4'd3)&(w299|w271))
	                        |((I_t == 4'd4)&(w304|w296|w305|w279|w297))
	                        |((I_t == 4'd6)&(w306)));
	
	assign O_control[ 35] = (((I_t == 4'd5)&(w301|w302|w089|w050))
	                        |((I_t == 4'd3)&(w307|w075|w076))
	                        |((I_t == 4'd4)&(w308|w309|w083))
	                        |((I_t == 4'd2)&(w222|w095))
	                        |((I_t == 4'd6)&(w306))
	                        |((I_t == 4'd1)&(w096)));
	
	assign O_control[ 36] = (((I_t == 4'd3)&(w310|w004|w033|w017)));
	
	assign O_control[ 37] = (((I_t == 4'd1)&(w311)));
	
	assign O_control[ 38] = (((I_t == 4'd1)&(w312)));
	
	assign O_control[ 39] = (((I_t == 4'd1)&(w312)));
	
	assign O_control[ 40] = (((I_t == 4'd2)&(w000|w166|w002|w313|w169|w038|w006))
	                        |((I_t == 4'd3)&(w115|w116|w117|w118))
	                        |((I_t == 4'd1)&(w312)));
	
	assign O_control[ 41] = (((I_t == 4'd1)&(w312)));
	
	assign O_control[ 42] = (((I_t == 4'd1)&(w312)));
	
	assign O_control[ 43] = (((I_t == 4'd3)&(w110|w047|w041|w163|w043|w006))
	                        |((I_t == 4'd4)&(w115|w116|w117|w118))
	                        |((I_t == 4'd2)&(w312)));
	
	assign O_control[ 44] = (((I_t == 4'd2)&(w312)));
	
	assign O_control[ 45] = (((I_t == 4'd3)&(w110|w047|w041|w163|w043|w006))
	                        |((I_t == 4'd4)&(w115|w116|w117|w118))
	                        |((I_t == 4'd2)&(w312)));
	
	assign O_control[ 46] = (((I_t == 4'd3)&(w312))
	                        |((I_t == 4'd2)&(w312)));
	
	assign O_control[ 47] = (((I_t == 4'd2)&(w312)));
	
	assign O_control[ 48] = (((I_t == 4'd2)&(w103|w314|w107|w038|w315)));
	
	assign O_control[ 49] = (((I_t == 4'd2)&(w115|w116|w117|w118)));
	
	assign O_control[ 50] = (((I_t == 4'd3)&(w115|w116|w117|w118))
	                        |((I_t == 4'd2)&(w316|w317|w318|w319|w320)));
	
	assign O_control[ 51] = (((I_t == 4'd2)&(w110|w321|w144|w235|w322|w163|w323))
	                        |((I_t == 4'd3)&(w115|w117|w179)));
	
	assign O_control[ 52] = (((I_t == 4'd1)&(w324)));
	
	assign O_control[ 53] = (((I_t == 4'd4)&(w325|w211))
	                        |((I_t == 4'd5)&(w326|w327|w198|w328))
	                        |((I_t == 4'd7)&(w329))
	                        |((I_t == 4'd3)&(w330|w331|w332|w333))
	                        |((I_t == 4'd1)&(w334|w096))
	                        |((I_t == 4'd6)&(w335))
	                        |((I_t == 4'd2)&(w336|w337)));
	
	assign O_control[ 54] = (((I_t == 4'd4)&(w338|w339|w335))
	                        |((I_t == 4'd5)&(w300|w329))
	                        |((I_t == 4'd3)&(w340|w326|w327))
	                        |((I_t == 4'd2)&(w325))
	                        |((I_t == 4'd1)&(w341)));
	
	assign O_control[ 55] = (((I_t == 4'd2)&(w342))
	                        |((I_t == 4'd3)&(w343)));
	
	assign O_control[ 56] = (((I_t == 4'd2)&(w344|w069))
	                        |((I_t == 4'd4)&(w072))
	                        |((I_t == 4'd3)&(w344)));
	
	assign O_control[ 57] = (((I_t == 4'd3)&(w345|w072)));
	
	assign O_control[ 58] = (((I_t == 4'd1)&(w346)));
	
	assign O_control[ 59] = (((I_t == 4'd1)&(w347)));
	
	assign O_control[ 60] = (((I_t == 4'd4)&(w072))
	                        |((I_t == 4'd3)&(w162)));
	
	assign O_control[ 61] = (((I_t == 4'd5)&(w072))
	                        |((I_t == 4'd4)&(w162)));
	
	assign O_control[ 62] = (((I_t == 4'd5)&(w348|w349|w350))
	                        |((I_t == 4'd1)&(w351))
	                        |((I_t == 4'd4)&(w352|w353))
	                        |((I_t == 4'd3)&(w354|w355))
	                        |((I_t == 4'd7)&(w356))
	                        |((I_t == 4'd2)&(w357))
	                        |((I_t == 4'd6)&(w358)));
	
	assign O_control[ 63] = (((I_t == 4'd3)&(w359|w348|w349))
	                        |((I_t == 4'd5)&(w360|w356|w361))
	                        |((I_t == 4'd4)&(w362|w358|w363))
	                        |((I_t == 4'd2)&(w352))
	                        |((I_t == 4'd1)&(w364))
	                        |((I_t == 4'd6)&(w365)));
	
	assign O_control[ 64] = (((I_t == 4'd1)&(w366)));
	
	assign O_control[ 65] = (((I_t == 4'd1)&(w367)));
	
	assign O_control[ 66] = (((I_t == 4'd3)&(w368|w369))
	                        |((I_t == 4'd5)&(w370|w371|w372))
	                        |((I_t == 4'd2)&(w373))
	                        |((I_t == 4'd4)&(w374|w375))
	                        |((I_t == 4'd6)&(w376))
	                        |((I_t == 4'd7)&(w377))
	                        |((I_t == 4'd1)&(w378)));
	
	assign O_control[ 67] = (((I_t == 4'd3)&(w379|w370|w371))
	                        |((I_t == 4'd4)&(w380|w381|w376))
	                        |((I_t == 4'd1)&(w382))
	                        |((I_t == 4'd5)&(w383|w377))
	                        |((I_t == 4'd2)&(w374)));
	
	assign O_control[ 68] = (((I_t == 4'd3)&(w229|w231|w232))
	                        |((I_t == 4'd2)&(w240))
	                        |((I_t == 4'd1)&(w236|w149))
	                        |((I_t == 4'd4)&(w144|w384))
	                        |((I_t == 4'd5)&(w057)));
	
	assign O_control[ 69] = (((I_t == 4'd2)&(w109)));
	
	assign O_control[ 70] = (((I_t == 4'd1)&(w385)));
	
	assign O_control[ 71] = (((I_t == 4'd1)&(w386)));
	
	assign O_control[ 72] = (((I_t == 4'd3)&(w332|w333))
	                        |((I_t == 4'd5)&(w328))
	                        |((I_t == 4'd1)&(w096))
	                        |((I_t == 4'd2)&(w337)));
	
	assign O_control[ 73] = (((I_t == 4'd3)&(w332|w333))
	                        |((I_t == 4'd5)&(w328))
	                        |((I_t == 4'd1)&(w096))
	                        |((I_t == 4'd2)&(w337)));
	
	assign O_control[ 74] = (((I_t == 4'd3)&(w387|w388))
	                        |((I_t == 4'd1)&(w389|w390|w391))
	                        |((I_t == 4'd2)&(w392)));
	
	assign O_control[ 75] = (((I_t == 4'd2)&(w393|w394))
	                        |((I_t == 4'd3)&(w395|w396|w397))
	                        |((I_t == 4'd1)&(w398|w399)));
	
	assign O_control[ 76] = (((I_t == 4'd5)&(w400|w401))
	                        |((I_t == 4'd2)&(w402))
	                        |((I_t == 4'd4)&(w403|w404|w405))
	                        |((I_t == 4'd3)&(w406|w407|w408))
	                        |((I_t == 4'd1)&(w409|w410)));
	
	assign O_control[ 77] = (((I_t == 4'd2)&(w411))
	                        |((I_t == 4'd1)&(w412|w391))
	                        |((I_t == 4'd3)&(w413|w414))
	                        |((I_t == 4'd4)&(w415)));
	
	assign O_control[ 78] = (((I_t == 4'd1)&(w256|w219|w416|w417)));
	
	assign O_control[ 79] = (((I_t == 4'd1)&(w418)));
	
	assign O_control[ 80] = (((I_t == 4'd1)&(w419)));
	
	assign O_control[ 81] = (((I_t == 4'd1)&(w420|w421|w416|w410|w422))
	                        |((I_t == 4'd3)&(w423|w424))
	                        |((I_t == 4'd4)&(w425))
	                        |((I_t == 4'd2)&(w426))
	                        |((I_t == 4'd5)&(w427)));
	
	assign O_control[ 82] = (((I_t == 4'd1)&(w428)));
	
	assign O_control[ 83] = (((I_t == 4'd1)&(w429)));
	
	assign O_control[ 84] = (((I_t == 4'd1)&(w430)));
	
	assign O_control[ 85] = (((I_t == 4'd2)&(w431|w432))
	                        |((I_t == 4'd3)&(w402|w433|w434|w435))
	                        |((I_t == 4'd4)&(w407|w408|w436))
	                        |((I_t == 4'd1)&(w437|w237))
	                        |((I_t == 4'd5)&(w405|w438))
	                        |((I_t == 4'd6)&(w401)));
	
	assign O_control[ 86] = (((I_t == 4'd3)&(w207))
	                        |((I_t == 4'd4)&(w213|w214))
	                        |((I_t == 4'd5)&(w002))
	                        |((I_t == 4'd6)&(w093)));
	
	assign O_control[ 87] = (((I_t == 4'd4)&(w439|w440|w245))
	                        |((I_t == 4'd3)&(w441|w252|w253))
	                        |((I_t == 4'd5)&(w442|w255))
	                        |((I_t == 4'd1)&(w443))
	                        |((I_t == 4'd2)&(w248)));
	
	assign O_control[ 88] = (((I_t == 4'd1)&(w444)));
	
	assign O_control[ 89] = (((I_t == 4'd1)&(w445)));
	
	assign O_control[ 90] = (((I_t == 4'd3)&(w248|w446|w447))
	                        |((I_t == 4'd5)&(w245|w448))
	                        |((I_t == 4'd6)&(w255))
	                        |((I_t == 4'd4)&(w252|w253|w449))
	                        |((I_t == 4'd1)&(w450))
	                        |((I_t == 4'd2)&(w451)));
	
	assign O_control[ 91] = (((I_t == 4'd1)&(w452)));
	
	assign O_control[ 92] = (((I_t == 4'd1)&(w453)));
	
	assign O_control[ 93] = (((I_t == 4'd0)));
	
	assign O_control[ 94] = (((I_t == 4'd0)));
	
endmodule