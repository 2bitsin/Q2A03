
	if (((curr_cycle == 2)&((curr_ir == 8'h5F)|(curr_ir == 8'h8F)|(curr_ir == 8'h4E)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'h2C)|(curr_ir == 8'hED)|(curr_ir == 8'hDD)|(curr_ir == 8'h79)|(curr_ir == 8'hDC)|(curr_ir == 8'h8D)|(curr_ir == 8'h2F)|(curr_ir == 8'h7C)|(curr_ir == 8'h1E)|(curr_ir == 8'hDF)|(curr_ir == 8'hFF)|(curr_ir == 8'h4F)|(curr_ir == 8'hCC)|(curr_ir == 8'hDE)|(curr_ir == 8'hCE)|(curr_ir == 8'h19)|(curr_ir == 8'h8E)|(curr_ir == 8'h99)|(curr_ir == 8'h3E)|(curr_ir == 8'h2E)|(curr_ir == 8'h7E)|(curr_ir == 8'h6E)|(curr_ir == 8'hCD)|(curr_ir == 8'h39)|(curr_ir == 8'h2D)|(curr_ir == 8'hBE)|(curr_ir == 8'h1C)|(curr_ir == 8'h7D)|(curr_ir == 8'hF9)|(curr_ir == 8'hBD)|(curr_ir == 8'hAD)|(curr_ir == 8'h6C)|(curr_ir == 8'hAC)|(curr_ir == 8'h1D)|(curr_ir == 8'h5D)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h0C)|(curr_ir == 8'h4C)|(curr_ir == 8'h1F)|(curr_ir == 8'hFC)|(curr_ir == 8'h6F)|(curr_ir == 8'hBC)|(curr_ir == 8'h5E)|(curr_ir == 8'h0E)|(curr_ir == 8'hDB)|(curr_ir == 8'hCF)|(curr_ir == 8'hFB)|(curr_ir == 8'h5B)|(curr_ir == 8'hFD)|(curr_ir == 8'h6D)|(curr_ir == 8'hEC)|(curr_ir == 8'h5C)|(curr_ir == 8'hD9)|(curr_ir == 8'h0D)|(curr_ir == 8'h4D)|(curr_ir == 8'hAE)|(curr_ir == 8'hB9)|(curr_ir == 8'h9D)|(curr_ir == 8'h8C)|(curr_ir == 8'hEF)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h3C)|(curr_ir == 8'hBF)|(curr_ir == 8'hAF)|(curr_ir == 8'h1B)|(curr_ir == 8'h0F)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h5A)|(curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'hC3)|(curr_ir == 8'h65)|(curr_ir == 8'hCD)|(curr_ir == 8'h49)|(curr_ir == 8'h8E)|(curr_ir == 8'hCE)|(curr_ir == 8'hB2)|(curr_ir == 8'hA2)|(curr_ir == 8'h2E)|(curr_ir == 8'h7D)|(curr_ir == 8'hBD)|(curr_ir == 8'h25)|(curr_ir == 8'hA1)|(curr_ir == 8'h09)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'h2D)|(curr_ir == 8'h6C)|(curr_ir == 8'hAC)|(curr_ir == 8'h90)|(curr_ir == 8'hF1)|(curr_ir == 8'h5D)|(curr_ir == 8'h38)|(curr_ir == 8'hD5)|(curr_ir == 8'h41)|(curr_ir == 8'h1C)|(curr_ir == 8'h05)|(curr_ir == 8'hE0)|(curr_ir == 8'h4C)|(curr_ir == 8'hC4)|(curr_ir == 8'h40)|(curr_ir == 8'h30)|(curr_ir == 8'h91)|(curr_ir == 8'h75)|(curr_ir == 8'hB5)|(curr_ir == 8'h1D)|(curr_ir == 8'h80)|(curr_ir == 8'h74)|(curr_ir == 8'h64)|(curr_ir == 8'hA4)|(curr_ir == 8'h0C)|(curr_ir == 8'hE9)|(curr_ir == 8'h7F)|(curr_ir == 8'h6F)|(curr_ir == 8'h63)|(curr_ir == 8'hF4)|(curr_ir == 8'hE8)|(curr_ir == 8'hD8)|(curr_ir == 8'hBC)|(curr_ir == 8'hFC)|(curr_ir == 8'h52)|(curr_ir == 8'hB3)|(curr_ir == 8'hF3)|(curr_ir == 8'hE3)|(curr_ir == 8'hD7)|(curr_ir == 8'hC7)|(curr_ir == 8'h3F)|(curr_ir == 8'h88)|(curr_ir == 8'h86)|(curr_ir == 8'h14)|(curr_ir == 8'hC6)|(curr_ir == 8'h53)|(curr_ir == 8'hFB)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h5B)|(curr_ir == 8'h1F)|(curr_ir == 8'h0F)|(curr_ir == 8'h03)|(curr_ir == 8'hFA)|(curr_ir == 8'h66)|(curr_ir == 8'h4A)|(curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'hAB)|(curr_ir == 8'hEB)|(curr_ir == 8'hDB)|(curr_ir == 8'hCF)|(curr_ir == 8'h55)|(curr_ir == 8'hB6)|(curr_ir == 8'h9A)|(curr_ir == 8'h06)|(curr_ir == 8'hDA)|(curr_ir == 8'h42)|(curr_ir == 8'hBE)|(curr_ir == 8'h26)|(curr_ir == 8'hA5)|(curr_ir == 8'h99)|(curr_ir == 8'h89)|(curr_ir == 8'h6D)|(curr_ir == 8'hEA)|(curr_ir == 8'h31)|(curr_ir == 8'h3A)|(curr_ir == 8'h15)|(curr_ir == 8'h7A)|(curr_ir == 8'hF2)|(curr_ir == 8'hD9)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'hE1)|(curr_ir == 8'h4D)|(curr_ir == 8'hAE)|(curr_ir == 8'h44)|(curr_ir == 8'hEC)|(curr_ir == 8'hB9)|(curr_ir == 8'hAD)|(curr_ir == 8'h9D)|(curr_ir == 8'h81)|(curr_ir == 8'hC1)|(curr_ir == 8'hE2)|(curr_ir == 8'h29)|(curr_ir == 8'h0D)|(curr_ir == 8'h78)|(curr_ir == 8'h5C)|(curr_ir == 8'hA8)|(curr_ir == 8'h8C)|(curr_ir == 8'h04)|(curr_ir == 8'hD1)|(curr_ir == 8'h28)|(curr_ir == 8'h18)|(curr_ir == 8'hF5)|(curr_ir == 8'hD0)|(curr_ir == 8'hC0)|(curr_ir == 8'h3C)|(curr_ir == 8'h17)|(curr_ir == 8'hB4)|(curr_ir == 8'h20)|(curr_ir == 8'hBF)|(curr_ir == 8'hA3)|(curr_ir == 8'h70)|(curr_ir == 8'h54)|(curr_ir == 8'h94)|(curr_ir == 8'h1A)|(curr_ir == 8'h92)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'h07)|(curr_ir == 8'h83)|(curr_ir == 8'hE4)|(curr_ir == 8'hC8)|(curr_ir == 8'h6A)|(curr_ir == 8'h5E)|(curr_ir == 8'h4E)|(curr_ir == 8'h12)|(curr_ir == 8'hEF)|(curr_ir == 8'hD3)|(curr_ir == 8'h3B)|(curr_ir == 8'hB7)|(curr_ir == 8'h59)|(curr_ir == 8'h82)|(curr_ir == 8'hDE)|(curr_ir == 8'hD2)|(curr_ir == 8'hC2)|(curr_ir == 8'h2A)|(curr_ir == 8'hA6)|(curr_ir == 8'h32)|(curr_ir == 8'h71)|(curr_ir == 8'hB1)|(curr_ir == 8'h19)|(curr_ir == 8'hF6)|(curr_ir == 8'h72)|(curr_ir == 8'h62)|(curr_ir == 8'h56)|(curr_ir == 8'h0A)|(curr_ir == 8'hA7)|(curr_ir == 8'hE7)|(curr_ir == 8'hE5)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h45)|(curr_ir == 8'h96)|(curr_ir == 8'h8A)|(curr_ir == 8'hD6)|(curr_ir == 8'hCA)|(curr_ir == 8'hBA)|(curr_ir == 8'h22)|(curr_ir == 8'h50)|(curr_ir == 8'h34)|(curr_ir == 8'h95)|(curr_ir == 8'h85)|(curr_ir == 8'h01)|(curr_ir == 8'h79)|(curr_ir == 8'hC5)|(curr_ir == 8'h3D)|(curr_ir == 8'h21)|(curr_ir == 8'h11)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'hA0)|(curr_ir == 8'h84)|(curr_ir == 8'h68)|(curr_ir == 8'h2C)|(curr_ir == 8'hC9)|(curr_ir == 8'h35)|(curr_ir == 8'h10)|(curr_ir == 8'hF9)|(curr_ir == 8'hED)|(curr_ir == 8'hDD)|(curr_ir == 8'h73)|(curr_ir == 8'h57)|(curr_ir == 8'hB8)|(curr_ir == 8'hF8)|(curr_ir == 8'hDC)|(curr_ir == 8'h48)|(curr_ir == 8'h69)|(curr_ir == 8'hA9)|(curr_ir == 8'h8D)|(curr_ir == 8'h2F)|(curr_ir == 8'hCB)|(curr_ir == 8'h37)|(curr_ir == 8'h58)|(curr_ir == 8'h98)|(curr_ir == 8'h00)|(curr_ir == 8'h7C)|(curr_ir == 8'h60)|(curr_ir == 8'h24)|(curr_ir == 8'h08)|(curr_ir == 8'h97)|(curr_ir == 8'h87)|(curr_ir == 8'hFF)|(curr_ir == 8'hCC)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'hB0)|(curr_ir == 8'hF0)|(curr_ir == 8'hD4)|(curr_ir == 8'h76)|(curr_ir == 8'h1E)|(curr_ir == 8'h27)|(curr_ir == 8'h02)|(curr_ir == 8'hAF)|(curr_ir == 8'h1B)|(curr_ir == 8'hDF)|(curr_ir == 8'h47)|(curr_ir == 8'hAA)|(curr_ir == 8'h16)|(curr_ir == 8'h46)|(curr_ir == 8'h36)|(curr_ir == 8'h4F)|(curr_ir == 8'h8F)|(curr_ir == 8'hF7)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h60)|(curr_ir == 8'h20)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hD0)|(curr_ir == 8'h70)|(curr_ir == 8'h50)|(curr_ir == 8'h10)|(curr_ir == 8'hB0)|(curr_ir == 8'hF0)|(curr_ir == 8'h90)|(curr_ir == 8'h30)))|
	    ((curr_cycle == 0)))
		G_addr = curr_pc;
	
	if (((curr_cycle == 2)&((curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'h8F)|(curr_ir == 8'h83)|(curr_ir == 8'h4E)|(curr_ir == 8'hC3)|(curr_ir == 8'hB7)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'h21)|(curr_ir == 8'hFE)|(curr_ir == 8'hE7)|(curr_ir == 8'hA6)|(curr_ir == 8'h71)|(curr_ir == 8'hD6)|(curr_ir == 8'hB1)|(curr_ir == 8'h95)|(curr_ir == 8'hF6)|(curr_ir == 8'hA7)|(curr_ir == 8'hC5)|(curr_ir == 8'h11)|(curr_ir == 8'hE5)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'hEE)|(curr_ir == 8'h35)|(curr_ir == 8'h96)|(curr_ir == 8'h2C)|(curr_ir == 8'h10)|(curr_ir == 8'h50)|(curr_ir == 8'h40)|(curr_ir == 8'hED)|(curr_ir == 8'hDD)|(curr_ir == 8'h01)|(curr_ir == 8'h79)|(curr_ir == 8'h74)|(curr_ir == 8'h68)|(curr_ir == 8'h73)|(curr_ir == 8'h57)|(curr_ir == 8'h24)|(curr_ir == 8'hDC)|(curr_ir == 8'h8D)|(curr_ir == 8'h46)|(curr_ir == 8'h2F)|(curr_ir == 8'h13)|(curr_ir == 8'hF0)|(curr_ir == 8'h37)|(curr_ir == 8'hD4)|(curr_ir == 8'h7C)|(curr_ir == 8'h1E)|(curr_ir == 8'h60)|(curr_ir == 8'hDF)|(curr_ir == 8'h47)|(curr_ir == 8'hFF)|(curr_ir == 8'h4F)|(curr_ir == 8'hCC)|(curr_ir == 8'hB0)|(curr_ir == 8'hDE)|(curr_ir == 8'hCE)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'hF7)|(curr_ir == 8'h27)|(curr_ir == 8'h25)|(curr_ir == 8'h19)|(curr_ir == 8'h65)|(curr_ir == 8'h16)|(curr_ir == 8'h8E)|(curr_ir == 8'h99)|(curr_ir == 8'h05)|(curr_ir == 8'h3E)|(curr_ir == 8'h2E)|(curr_ir == 8'h7E)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'hCD)|(curr_ir == 8'h39)|(curr_ir == 8'h2D)|(curr_ir == 8'hBE)|(curr_ir == 8'hF1)|(curr_ir == 8'h1C)|(curr_ir == 8'h7D)|(curr_ir == 8'hF9)|(curr_ir == 8'hBD)|(curr_ir == 8'hAD)|(curr_ir == 8'hA1)|(curr_ir == 8'h91)|(curr_ir == 8'h6C)|(curr_ir == 8'hAC)|(curr_ir == 8'hB5)|(curr_ir == 8'h90)|(curr_ir == 8'h1D)|(curr_ir == 8'h5D)|(curr_ir == 8'hD5)|(curr_ir == 8'h41)|(curr_ir == 8'hF3)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h0C)|(curr_ir == 8'h4C)|(curr_ir == 8'hC4)|(curr_ir == 8'h30)|(curr_ir == 8'h14)|(curr_ir == 8'h75)|(curr_ir == 8'hB3)|(curr_ir == 8'h1F)|(curr_ir == 8'hFC)|(curr_ir == 8'h64)|(curr_ir == 8'hA4)|(curr_ir == 8'h6F)|(curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'hBC)|(curr_ir == 8'h5E)|(curr_ir == 8'h03)|(curr_ir == 8'hD7)|(curr_ir == 8'hC7)|(curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'hC6)|(curr_ir == 8'hDB)|(curr_ir == 8'hCF)|(curr_ir == 8'hFB)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h5B)|(curr_ir == 8'h26)|(curr_ir == 8'h66)|(curr_ir == 8'h56)|(curr_ir == 8'h31)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'hB6)|(curr_ir == 8'h06)|(curr_ir == 8'h04)|(curr_ir == 8'hFD)|(curr_ir == 8'h44)|(curr_ir == 8'hA5)|(curr_ir == 8'h6D)|(curr_ir == 8'hEC)|(curr_ir == 8'h5C)|(curr_ir == 8'hD9)|(curr_ir == 8'h45)|(curr_ir == 8'hC1)|(curr_ir == 8'h0D)|(curr_ir == 8'hE1)|(curr_ir == 8'h4D)|(curr_ir == 8'hAE)|(curr_ir == 8'h34)|(curr_ir == 8'h28)|(curr_ir == 8'hD0)|(curr_ir == 8'hF5)|(curr_ir == 8'hB9)|(curr_ir == 8'h9D)|(curr_ir == 8'h81)|(curr_ir == 8'h23)|(curr_ir == 8'h17)|(curr_ir == 8'hF4)|(curr_ir == 8'hE4)|(curr_ir == 8'h8C)|(curr_ir == 8'h70)|(curr_ir == 8'hD1)|(curr_ir == 8'hEF)|(curr_ir == 8'hE3)|(curr_ir == 8'h3B)|(curr_ir == 8'h97)|(curr_ir == 8'h7B)|(curr_ir == 8'h3C)|(curr_ir == 8'hB4)|(curr_ir == 8'h20)|(curr_ir == 8'h07)|(curr_ir == 8'hBF)|(curr_ir == 8'hAF)|(curr_ir == 8'h1B)|(curr_ir == 8'hA3)|(curr_ir == 8'h0F)|(curr_ir == 8'h54)|(curr_ir == 8'h94)|(curr_ir == 8'hD3)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h5A)|(curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'hC3)|(curr_ir == 8'h65)|(curr_ir == 8'hCD)|(curr_ir == 8'h49)|(curr_ir == 8'h8E)|(curr_ir == 8'hCE)|(curr_ir == 8'hB2)|(curr_ir == 8'hA2)|(curr_ir == 8'h2E)|(curr_ir == 8'h7D)|(curr_ir == 8'hBD)|(curr_ir == 8'h25)|(curr_ir == 8'hA1)|(curr_ir == 8'h09)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'h2D)|(curr_ir == 8'h6C)|(curr_ir == 8'hAC)|(curr_ir == 8'h90)|(curr_ir == 8'hF1)|(curr_ir == 8'h5D)|(curr_ir == 8'h38)|(curr_ir == 8'hD5)|(curr_ir == 8'h41)|(curr_ir == 8'h1C)|(curr_ir == 8'h05)|(curr_ir == 8'hE0)|(curr_ir == 8'h4C)|(curr_ir == 8'hC4)|(curr_ir == 8'h40)|(curr_ir == 8'h30)|(curr_ir == 8'h91)|(curr_ir == 8'h75)|(curr_ir == 8'hB5)|(curr_ir == 8'h1D)|(curr_ir == 8'h80)|(curr_ir == 8'h74)|(curr_ir == 8'h64)|(curr_ir == 8'hA4)|(curr_ir == 8'h0C)|(curr_ir == 8'hE9)|(curr_ir == 8'h7F)|(curr_ir == 8'h6F)|(curr_ir == 8'h63)|(curr_ir == 8'hF4)|(curr_ir == 8'hE8)|(curr_ir == 8'hD8)|(curr_ir == 8'hBC)|(curr_ir == 8'hFC)|(curr_ir == 8'h52)|(curr_ir == 8'hB3)|(curr_ir == 8'hF3)|(curr_ir == 8'hE3)|(curr_ir == 8'hD7)|(curr_ir == 8'hC7)|(curr_ir == 8'h3F)|(curr_ir == 8'h88)|(curr_ir == 8'h86)|(curr_ir == 8'h14)|(curr_ir == 8'hC6)|(curr_ir == 8'h53)|(curr_ir == 8'hFB)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h5B)|(curr_ir == 8'h1F)|(curr_ir == 8'h0F)|(curr_ir == 8'h03)|(curr_ir == 8'hFA)|(curr_ir == 8'h66)|(curr_ir == 8'h4A)|(curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'hAB)|(curr_ir == 8'hEB)|(curr_ir == 8'hDB)|(curr_ir == 8'hCF)|(curr_ir == 8'h55)|(curr_ir == 8'hB6)|(curr_ir == 8'h9A)|(curr_ir == 8'h06)|(curr_ir == 8'hDA)|(curr_ir == 8'h42)|(curr_ir == 8'hBE)|(curr_ir == 8'h26)|(curr_ir == 8'hA5)|(curr_ir == 8'h99)|(curr_ir == 8'h89)|(curr_ir == 8'h6D)|(curr_ir == 8'hEA)|(curr_ir == 8'h31)|(curr_ir == 8'h3A)|(curr_ir == 8'h15)|(curr_ir == 8'h7A)|(curr_ir == 8'hF2)|(curr_ir == 8'hD9)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'hE1)|(curr_ir == 8'h4D)|(curr_ir == 8'hAE)|(curr_ir == 8'h44)|(curr_ir == 8'hEC)|(curr_ir == 8'hB9)|(curr_ir == 8'hAD)|(curr_ir == 8'h9D)|(curr_ir == 8'h81)|(curr_ir == 8'hC1)|(curr_ir == 8'hE2)|(curr_ir == 8'h29)|(curr_ir == 8'h0D)|(curr_ir == 8'h78)|(curr_ir == 8'h5C)|(curr_ir == 8'hA8)|(curr_ir == 8'h8C)|(curr_ir == 8'h04)|(curr_ir == 8'hD1)|(curr_ir == 8'h28)|(curr_ir == 8'h18)|(curr_ir == 8'hF5)|(curr_ir == 8'hD0)|(curr_ir == 8'hC0)|(curr_ir == 8'h3C)|(curr_ir == 8'h17)|(curr_ir == 8'hB4)|(curr_ir == 8'h20)|(curr_ir == 8'hBF)|(curr_ir == 8'hA3)|(curr_ir == 8'h70)|(curr_ir == 8'h54)|(curr_ir == 8'h94)|(curr_ir == 8'h1A)|(curr_ir == 8'h92)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'h07)|(curr_ir == 8'h83)|(curr_ir == 8'hE4)|(curr_ir == 8'hC8)|(curr_ir == 8'h6A)|(curr_ir == 8'h5E)|(curr_ir == 8'h4E)|(curr_ir == 8'h12)|(curr_ir == 8'hEF)|(curr_ir == 8'hD3)|(curr_ir == 8'h3B)|(curr_ir == 8'hB7)|(curr_ir == 8'h59)|(curr_ir == 8'h82)|(curr_ir == 8'hDE)|(curr_ir == 8'hD2)|(curr_ir == 8'hC2)|(curr_ir == 8'h2A)|(curr_ir == 8'hA6)|(curr_ir == 8'h32)|(curr_ir == 8'h71)|(curr_ir == 8'hB1)|(curr_ir == 8'h19)|(curr_ir == 8'hF6)|(curr_ir == 8'h72)|(curr_ir == 8'h62)|(curr_ir == 8'h56)|(curr_ir == 8'h0A)|(curr_ir == 8'hA7)|(curr_ir == 8'hE7)|(curr_ir == 8'hE5)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h45)|(curr_ir == 8'h96)|(curr_ir == 8'h8A)|(curr_ir == 8'hD6)|(curr_ir == 8'hBA)|(curr_ir == 8'hCA)|(curr_ir == 8'h22)|(curr_ir == 8'h50)|(curr_ir == 8'h34)|(curr_ir == 8'h95)|(curr_ir == 8'h85)|(curr_ir == 8'h01)|(curr_ir == 8'h79)|(curr_ir == 8'hC5)|(curr_ir == 8'h3D)|(curr_ir == 8'h21)|(curr_ir == 8'h11)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'hA0)|(curr_ir == 8'h84)|(curr_ir == 8'h68)|(curr_ir == 8'h2C)|(curr_ir == 8'hC9)|(curr_ir == 8'h35)|(curr_ir == 8'h10)|(curr_ir == 8'hF9)|(curr_ir == 8'hED)|(curr_ir == 8'hDD)|(curr_ir == 8'h73)|(curr_ir == 8'h57)|(curr_ir == 8'hB8)|(curr_ir == 8'hF8)|(curr_ir == 8'hDC)|(curr_ir == 8'h48)|(curr_ir == 8'h69)|(curr_ir == 8'hA9)|(curr_ir == 8'h8D)|(curr_ir == 8'h2F)|(curr_ir == 8'h37)|(curr_ir == 8'h58)|(curr_ir == 8'h98)|(curr_ir == 8'h00)|(curr_ir == 8'h7C)|(curr_ir == 8'h60)|(curr_ir == 8'h24)|(curr_ir == 8'h08)|(curr_ir == 8'h97)|(curr_ir == 8'h87)|(curr_ir == 8'hFF)|(curr_ir == 8'hCC)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'hB0)|(curr_ir == 8'hF0)|(curr_ir == 8'hD4)|(curr_ir == 8'h76)|(curr_ir == 8'h1E)|(curr_ir == 8'h02)|(curr_ir == 8'h27)|(curr_ir == 8'hAF)|(curr_ir == 8'h1B)|(curr_ir == 8'hDF)|(curr_ir == 8'h47)|(curr_ir == 8'hAA)|(curr_ir == 8'h16)|(curr_ir == 8'h46)|(curr_ir == 8'h36)|(curr_ir == 8'h4F)|(curr_ir == 8'h8F)|(curr_ir == 8'hF7)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'h53)|(curr_ir == 8'hB6)|(curr_ir == 8'h5E)|(curr_ir == 8'hFB)|(curr_ir == 8'h5B)|(curr_ir == 8'h56)|(curr_ir == 8'hDB)|(curr_ir == 8'hD9)|(curr_ir == 8'hCD)|(curr_ir == 8'hBE)|(curr_ir == 8'hAE)|(curr_ir == 8'hB9)|(curr_ir == 8'h31)|(curr_ir == 8'hAD)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'hFD)|(curr_ir == 8'hE1)|(curr_ir == 8'h4D)|(curr_ir == 8'h6D)|(curr_ir == 8'hEC)|(curr_ir == 8'hD0)|(curr_ir == 8'h3C)|(curr_ir == 8'h9D)|(curr_ir == 8'h81)|(curr_ir == 8'h5C)|(curr_ir == 8'hC1)|(curr_ir == 8'h0D)|(curr_ir == 8'h70)|(curr_ir == 8'h34)|(curr_ir == 8'hD1)|(curr_ir == 8'hF5)|(curr_ir == 8'h7B)|(curr_ir == 8'h6F)|(curr_ir == 8'h23)|(curr_ir == 8'h17)|(curr_ir == 8'hF4)|(curr_ir == 8'hBF)|(curr_ir == 8'hAF)|(curr_ir == 8'hA3)|(curr_ir == 8'hEF)|(curr_ir == 8'hD3)|(curr_ir == 8'hE3)|(curr_ir == 8'h3B)|(curr_ir == 8'h5F)|(curr_ir == 8'hDE)|(curr_ir == 8'h83)|(curr_ir == 8'h1B)|(curr_ir == 8'h0F)|(curr_ir == 8'h7E)|(curr_ir == 8'hB7)|(curr_ir == 8'h4F)|(curr_ir == 8'h43)|(curr_ir == 8'h61)|(curr_ir == 8'h4E)|(curr_ir == 8'h3E)|(curr_ir == 8'hB1)|(curr_ir == 8'h19)|(curr_ir == 8'h59)|(curr_ir == 8'h79)|(curr_ir == 8'hF6)|(curr_ir == 8'h3D)|(curr_ir == 8'h21)|(curr_ir == 8'hFE)|(curr_ir == 8'h51)|(curr_ir == 8'h2C)|(curr_ir == 8'h71)|(curr_ir == 8'hED)|(curr_ir == 8'hD6)|(curr_ir == 8'h01)|(curr_ir == 8'h50)|(curr_ir == 8'h11)|(curr_ir == 8'hEE)|(curr_ir == 8'h35)|(curr_ir == 8'h10)|(curr_ir == 8'h40)|(curr_ir == 8'hDD)|(curr_ir == 8'hDC)|(curr_ir == 8'hCC)|(curr_ir == 8'hB0)|(curr_ir == 8'h68)|(curr_ir == 8'h37)|(curr_ir == 8'h73)|(curr_ir == 8'h63)|(curr_ir == 8'h7C)|(curr_ir == 8'h57)|(curr_ir == 8'h60)|(curr_ir == 8'hFF)|(curr_ir == 8'h2F)|(curr_ir == 8'h13)|(curr_ir == 8'hF0)|(curr_ir == 8'hD4)|(curr_ir == 8'h76)|(curr_ir == 8'h1E)|(curr_ir == 8'hDF)|(curr_ir == 8'hCF)|(curr_ir == 8'hC3)|(curr_ir == 8'hCE)|(curr_ir == 8'h36)|(curr_ir == 8'hF7)|(curr_ir == 8'h99)|(curr_ir == 8'hBD)|(curr_ir == 8'h6E)|(curr_ir == 8'h16)|(curr_ir == 8'hF1)|(curr_ir == 8'h5D)|(curr_ir == 8'h7D)|(curr_ir == 8'h2E)|(curr_ir == 8'hA1)|(curr_ir == 8'h91)|(curr_ir == 8'h75)|(curr_ir == 8'h39)|(curr_ir == 8'h2D)|(curr_ir == 8'h1D)|(curr_ir == 8'hAC)|(curr_ir == 8'h90)|(curr_ir == 8'h74)|(curr_ir == 8'h28)|(curr_ir == 8'hD5)|(curr_ir == 8'h41)|(curr_ir == 8'h1C)|(curr_ir == 8'hF9)|(curr_ir == 8'h7F)|(curr_ir == 8'hB4)|(curr_ir == 8'h6C)|(curr_ir == 8'hB5)|(curr_ir == 8'hB3)|(curr_ir == 8'hF3)|(curr_ir == 8'hD7)|(curr_ir == 8'h3F)|(curr_ir == 8'h0C)|(curr_ir == 8'h30)|(curr_ir == 8'h14)|(curr_ir == 8'h77)|(curr_ir == 8'h1F)|(curr_ir == 8'hBC)|(curr_ir == 8'h03)|(curr_ir == 8'hFC)|(curr_ir == 8'h54)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h57)|(curr_ir == 8'h60)|(curr_ir == 8'hD3)|(curr_ir == 8'h43)|(curr_ir == 8'h71)|(curr_ir == 8'hB1)|(curr_ir == 8'h21)|(curr_ir == 8'h11)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h01)|(curr_ir == 8'h73)|(curr_ir == 8'h40)|(curr_ir == 8'h2F)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'h63)|(curr_ir == 8'h37)|(curr_ir == 8'hC3)|(curr_ir == 8'h4F)|(curr_ir == 8'hA1)|(curr_ir == 8'hF1)|(curr_ir == 8'h41)|(curr_ir == 8'h00)|(curr_ir == 8'hE3)|(curr_ir == 8'hF3)|(curr_ir == 8'h6F)|(curr_ir == 8'h20)|(curr_ir == 8'h77)|(curr_ir == 8'hB3)|(curr_ir == 8'hA3)|(curr_ir == 8'h0F)|(curr_ir == 8'h03)|(curr_ir == 8'h53)|(curr_ir == 8'h33)|(curr_ir == 8'h31)|(curr_ir == 8'hE1)|(curr_ir == 8'hC1)|(curr_ir == 8'hD1)|(curr_ir == 8'h17)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h1F)|(curr_ir == 8'h3F)|(curr_ir == 8'h5B)|(curr_ir == 8'h1B)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h00)|(curr_ir == 8'h7F)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h27)|(curr_ir == 8'h60)|(curr_ir == 8'hFF)|(curr_ir == 8'h5B)|(curr_ir == 8'h3E)|(curr_ir == 8'hDF)|(curr_ir == 8'hC3)|(curr_ir == 8'h7D)|(curr_ir == 8'hBD)|(curr_ir == 8'hA1)|(curr_ir == 8'h6C)|(curr_ir == 8'h1D)|(curr_ir == 8'hF1)|(curr_ir == 8'h11)|(curr_ir == 8'h5D)|(curr_ir == 8'h41)|(curr_ir == 8'h1C)|(curr_ir == 8'h91)|(curr_ir == 8'hF9)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h63)|(curr_ir == 8'hB3)|(curr_ir == 8'hA3)|(curr_ir == 8'h1F)|(curr_ir == 8'hF3)|(curr_ir == 8'h03)|(curr_ir == 8'hFC)|(curr_ir == 8'h1E)|(curr_ir == 8'h53)|(curr_ir == 8'hBC)|(curr_ir == 8'h5E)|(curr_ir == 8'hE3)|(curr_ir == 8'h33)|(curr_ir == 8'h31)|(curr_ir == 8'hFB)|(curr_ir == 8'h67)|(curr_ir == 8'hD9)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'hBE)|(curr_ir == 8'hB9)|(curr_ir == 8'h5C)|(curr_ir == 8'hE1)|(curr_ir == 8'hD1)|(curr_ir == 8'hDC)|(curr_ir == 8'h3C)|(curr_ir == 8'h81)|(curr_ir == 8'hC1)|(curr_ir == 8'h07)|(curr_ir == 8'hBF)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'h1B)|(curr_ir == 8'hD3)|(curr_ir == 8'hDE)|(curr_ir == 8'hDB)|(curr_ir == 8'h83)|(curr_ir == 8'h7E)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'h21)|(curr_ir == 8'h61)|(curr_ir == 8'h71)|(curr_ir == 8'hB1)|(curr_ir == 8'h19)|(curr_ir == 8'h01)|(curr_ir == 8'h79)|(curr_ir == 8'hFE)|(curr_ir == 8'h51)|(curr_ir == 8'h40)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'h7C)|(curr_ir == 8'hDD)|(curr_ir == 8'h73)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h73)|(curr_ir == 8'h63)|(curr_ir == 8'h13)|(curr_ir == 8'h03)|(curr_ir == 8'h53)|(curr_ir == 8'h33)|(curr_ir == 8'h23)|(curr_ir == 8'h43)))|
	    ((curr_cycle == 0)))
		G_rdwr = 1;
	
	if (((curr_cycle == 2)&((curr_ir == 8'h43)|(curr_ir == 8'h8F)|(curr_ir == 8'h83)|(curr_ir == 8'h4E)|(curr_ir == 8'hC3)|(curr_ir == 8'hB7)|(curr_ir == 8'h21)|(curr_ir == 8'hFE)|(curr_ir == 8'hE7)|(curr_ir == 8'h71)|(curr_ir == 8'hD6)|(curr_ir == 8'hB1)|(curr_ir == 8'h95)|(curr_ir == 8'hF6)|(curr_ir == 8'h11)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'hEE)|(curr_ir == 8'h35)|(curr_ir == 8'h96)|(curr_ir == 8'h2C)|(curr_ir == 8'h00)|(curr_ir == 8'h40)|(curr_ir == 8'hED)|(curr_ir == 8'h01)|(curr_ir == 8'h74)|(curr_ir == 8'h68)|(curr_ir == 8'h73)|(curr_ir == 8'h57)|(curr_ir == 8'h8D)|(curr_ir == 8'h46)|(curr_ir == 8'h2F)|(curr_ir == 8'h13)|(curr_ir == 8'h37)|(curr_ir == 8'hD4)|(curr_ir == 8'h1E)|(curr_ir == 8'h60)|(curr_ir == 8'h47)|(curr_ir == 8'h4F)|(curr_ir == 8'hCC)|(curr_ir == 8'hDE)|(curr_ir == 8'hCE)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'hF7)|(curr_ir == 8'h27)|(curr_ir == 8'h16)|(curr_ir == 8'h8E)|(curr_ir == 8'h99)|(curr_ir == 8'h3E)|(curr_ir == 8'h2E)|(curr_ir == 8'h7E)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'hCD)|(curr_ir == 8'h2D)|(curr_ir == 8'hF1)|(curr_ir == 8'hAD)|(curr_ir == 8'hA1)|(curr_ir == 8'h91)|(curr_ir == 8'h6C)|(curr_ir == 8'hAC)|(curr_ir == 8'hB5)|(curr_ir == 8'hD5)|(curr_ir == 8'h41)|(curr_ir == 8'hF3)|(curr_ir == 8'h0C)|(curr_ir == 8'h14)|(curr_ir == 8'h75)|(curr_ir == 8'hB3)|(curr_ir == 8'h6F)|(curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'h5E)|(curr_ir == 8'h03)|(curr_ir == 8'hD7)|(curr_ir == 8'hC7)|(curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'hC6)|(curr_ir == 8'hCF)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h26)|(curr_ir == 8'h66)|(curr_ir == 8'h56)|(curr_ir == 8'h31)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'hB6)|(curr_ir == 8'h06)|(curr_ir == 8'h6D)|(curr_ir == 8'hEC)|(curr_ir == 8'hC1)|(curr_ir == 8'h0D)|(curr_ir == 8'hE1)|(curr_ir == 8'h4D)|(curr_ir == 8'hAE)|(curr_ir == 8'h34)|(curr_ir == 8'h28)|(curr_ir == 8'hF5)|(curr_ir == 8'h9D)|(curr_ir == 8'h81)|(curr_ir == 8'h23)|(curr_ir == 8'h17)|(curr_ir == 8'hF4)|(curr_ir == 8'h8C)|(curr_ir == 8'hD1)|(curr_ir == 8'hEF)|(curr_ir == 8'hE3)|(curr_ir == 8'h97)|(curr_ir == 8'hB4)|(curr_ir == 8'h20)|(curr_ir == 8'h07)|(curr_ir == 8'hAF)|(curr_ir == 8'hA3)|(curr_ir == 8'h0F)|(curr_ir == 8'h54)|(curr_ir == 8'h94)|(curr_ir == 8'hD3)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'hC3)|(curr_ir == 8'h65)|(curr_ir == 8'hCD)|(curr_ir == 8'h8E)|(curr_ir == 8'hCE)|(curr_ir == 8'h2E)|(curr_ir == 8'h7D)|(curr_ir == 8'hBD)|(curr_ir == 8'h25)|(curr_ir == 8'hA1)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'h2D)|(curr_ir == 8'h6C)|(curr_ir == 8'hAC)|(curr_ir == 8'hF1)|(curr_ir == 8'h5D)|(curr_ir == 8'hD5)|(curr_ir == 8'h41)|(curr_ir == 8'h1C)|(curr_ir == 8'h05)|(curr_ir == 8'h4C)|(curr_ir == 8'hC4)|(curr_ir == 8'h40)|(curr_ir == 8'h91)|(curr_ir == 8'h75)|(curr_ir == 8'hB5)|(curr_ir == 8'h1D)|(curr_ir == 8'h74)|(curr_ir == 8'h64)|(curr_ir == 8'hA4)|(curr_ir == 8'h0C)|(curr_ir == 8'h7F)|(curr_ir == 8'h6F)|(curr_ir == 8'h63)|(curr_ir == 8'hF4)|(curr_ir == 8'hBC)|(curr_ir == 8'hFC)|(curr_ir == 8'hB3)|(curr_ir == 8'hF3)|(curr_ir == 8'hE3)|(curr_ir == 8'hD7)|(curr_ir == 8'hC7)|(curr_ir == 8'h3F)|(curr_ir == 8'h86)|(curr_ir == 8'h14)|(curr_ir == 8'hC6)|(curr_ir == 8'h53)|(curr_ir == 8'hFB)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h5B)|(curr_ir == 8'h1F)|(curr_ir == 8'h0F)|(curr_ir == 8'h03)|(curr_ir == 8'h66)|(curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'hDB)|(curr_ir == 8'hCF)|(curr_ir == 8'h55)|(curr_ir == 8'hB6)|(curr_ir == 8'h06)|(curr_ir == 8'hBE)|(curr_ir == 8'h26)|(curr_ir == 8'hA5)|(curr_ir == 8'h99)|(curr_ir == 8'h6D)|(curr_ir == 8'h31)|(curr_ir == 8'h15)|(curr_ir == 8'hD9)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'hE1)|(curr_ir == 8'h4D)|(curr_ir == 8'hAE)|(curr_ir == 8'h44)|(curr_ir == 8'hEC)|(curr_ir == 8'hB9)|(curr_ir == 8'hAD)|(curr_ir == 8'h9D)|(curr_ir == 8'h81)|(curr_ir == 8'hC1)|(curr_ir == 8'h0D)|(curr_ir == 8'h5C)|(curr_ir == 8'h8C)|(curr_ir == 8'h04)|(curr_ir == 8'hD1)|(curr_ir == 8'h28)|(curr_ir == 8'hF5)|(curr_ir == 8'h3C)|(curr_ir == 8'h17)|(curr_ir == 8'hB4)|(curr_ir == 8'h20)|(curr_ir == 8'hBF)|(curr_ir == 8'hA3)|(curr_ir == 8'h54)|(curr_ir == 8'h94)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'h07)|(curr_ir == 8'h83)|(curr_ir == 8'hE4)|(curr_ir == 8'h5E)|(curr_ir == 8'h4E)|(curr_ir == 8'hEF)|(curr_ir == 8'hD3)|(curr_ir == 8'h3B)|(curr_ir == 8'hB7)|(curr_ir == 8'h59)|(curr_ir == 8'hDE)|(curr_ir == 8'hA6)|(curr_ir == 8'h71)|(curr_ir == 8'hB1)|(curr_ir == 8'h19)|(curr_ir == 8'hF6)|(curr_ir == 8'h56)|(curr_ir == 8'hA7)|(curr_ir == 8'hE7)|(curr_ir == 8'hE5)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h45)|(curr_ir == 8'h96)|(curr_ir == 8'hD6)|(curr_ir == 8'h34)|(curr_ir == 8'h95)|(curr_ir == 8'h85)|(curr_ir == 8'h01)|(curr_ir == 8'h79)|(curr_ir == 8'hC5)|(curr_ir == 8'h3D)|(curr_ir == 8'h21)|(curr_ir == 8'h11)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'h84)|(curr_ir == 8'h68)|(curr_ir == 8'h2C)|(curr_ir == 8'h35)|(curr_ir == 8'hF9)|(curr_ir == 8'hED)|(curr_ir == 8'hDD)|(curr_ir == 8'h73)|(curr_ir == 8'h57)|(curr_ir == 8'hDC)|(curr_ir == 8'h48)|(curr_ir == 8'h8D)|(curr_ir == 8'h2F)|(curr_ir == 8'h37)|(curr_ir == 8'h00)|(curr_ir == 8'h7C)|(curr_ir == 8'h60)|(curr_ir == 8'h24)|(curr_ir == 8'h08)|(curr_ir == 8'h97)|(curr_ir == 8'h87)|(curr_ir == 8'hFF)|(curr_ir == 8'hCC)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'hD4)|(curr_ir == 8'h76)|(curr_ir == 8'h1E)|(curr_ir == 8'h27)|(curr_ir == 8'hAF)|(curr_ir == 8'h1B)|(curr_ir == 8'hDF)|(curr_ir == 8'h47)|(curr_ir == 8'h16)|(curr_ir == 8'h46)|(curr_ir == 8'h36)|(curr_ir == 8'h4F)|(curr_ir == 8'h8F)|(curr_ir == 8'hF7)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hC7)|(curr_ir == 8'h0E)|(curr_ir == 8'hC6)|(curr_ir == 8'h5E)|(curr_ir == 8'hFB)|(curr_ir == 8'h67)|(curr_ir == 8'h5B)|(curr_ir == 8'h66)|(curr_ir == 8'h56)|(curr_ir == 8'hDB)|(curr_ir == 8'hD9)|(curr_ir == 8'hBE)|(curr_ir == 8'h26)|(curr_ir == 8'hB9)|(curr_ir == 8'h06)|(curr_ir == 8'hFD)|(curr_ir == 8'hE1)|(curr_ir == 8'h3C)|(curr_ir == 8'h9D)|(curr_ir == 8'h81)|(curr_ir == 8'h5C)|(curr_ir == 8'hC1)|(curr_ir == 8'h7B)|(curr_ir == 8'h6F)|(curr_ir == 8'h23)|(curr_ir == 8'h17)|(curr_ir == 8'h07)|(curr_ir == 8'hBF)|(curr_ir == 8'hA3)|(curr_ir == 8'hEF)|(curr_ir == 8'hE3)|(curr_ir == 8'h3B)|(curr_ir == 8'h5F)|(curr_ir == 8'hDE)|(curr_ir == 8'h83)|(curr_ir == 8'h1B)|(curr_ir == 8'h0F)|(curr_ir == 8'h7E)|(curr_ir == 8'hE7)|(curr_ir == 8'h4F)|(curr_ir == 8'h43)|(curr_ir == 8'h61)|(curr_ir == 8'h4E)|(curr_ir == 8'h3E)|(curr_ir == 8'h19)|(curr_ir == 8'h59)|(curr_ir == 8'h79)|(curr_ir == 8'hF6)|(curr_ir == 8'h3D)|(curr_ir == 8'h21)|(curr_ir == 8'hFE)|(curr_ir == 8'hD6)|(curr_ir == 8'h01)|(curr_ir == 8'hEE)|(curr_ir == 8'h00)|(curr_ir == 8'h40)|(curr_ir == 8'hDD)|(curr_ir == 8'hDC)|(curr_ir == 8'h37)|(curr_ir == 8'h63)|(curr_ir == 8'h7C)|(curr_ir == 8'h57)|(curr_ir == 8'h60)|(curr_ir == 8'hFF)|(curr_ir == 8'h46)|(curr_ir == 8'h2F)|(curr_ir == 8'h76)|(curr_ir == 8'h1E)|(curr_ir == 8'hDF)|(curr_ir == 8'hCF)|(curr_ir == 8'h47)|(curr_ir == 8'hC3)|(curr_ir == 8'hCE)|(curr_ir == 8'h36)|(curr_ir == 8'hF7)|(curr_ir == 8'h99)|(curr_ir == 8'h27)|(curr_ir == 8'hBD)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'h16)|(curr_ir == 8'h5D)|(curr_ir == 8'h7D)|(curr_ir == 8'h2E)|(curr_ir == 8'hA1)|(curr_ir == 8'h91)|(curr_ir == 8'h39)|(curr_ir == 8'h1D)|(curr_ir == 8'h41)|(curr_ir == 8'h1C)|(curr_ir == 8'hF9)|(curr_ir == 8'h7F)|(curr_ir == 8'h6C)|(curr_ir == 8'hD7)|(curr_ir == 8'h3F)|(curr_ir == 8'h20)|(curr_ir == 8'h77)|(curr_ir == 8'h1F)|(curr_ir == 8'hBC)|(curr_ir == 8'h03)|(curr_ir == 8'hFC)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hD7)|(curr_ir == 8'h37)|(curr_ir == 8'h60)|(curr_ir == 8'hFF)|(curr_ir == 8'h5B)|(curr_ir == 8'h4F)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'h3E)|(curr_ir == 8'hDF)|(curr_ir == 8'hCF)|(curr_ir == 8'hC3)|(curr_ir == 8'h16)|(curr_ir == 8'hCE)|(curr_ir == 8'hF7)|(curr_ir == 8'hA1)|(curr_ir == 8'h2E)|(curr_ir == 8'h6E)|(curr_ir == 8'hF1)|(curr_ir == 8'h11)|(curr_ir == 8'h41)|(curr_ir == 8'h91)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h63)|(curr_ir == 8'hB3)|(curr_ir == 8'hA3)|(curr_ir == 8'h1F)|(curr_ir == 8'hF3)|(curr_ir == 8'h03)|(curr_ir == 8'h1E)|(curr_ir == 8'h0E)|(curr_ir == 8'h53)|(curr_ir == 8'h77)|(curr_ir == 8'h5E)|(curr_ir == 8'hE3)|(curr_ir == 8'h33)|(curr_ir == 8'h31)|(curr_ir == 8'hFB)|(curr_ir == 8'h56)|(curr_ir == 8'h17)|(curr_ir == 8'hE1)|(curr_ir == 8'hD1)|(curr_ir == 8'h20)|(curr_ir == 8'h81)|(curr_ir == 8'hC1)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h6F)|(curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'h1B)|(curr_ir == 8'hEF)|(curr_ir == 8'h0F)|(curr_ir == 8'hD3)|(curr_ir == 8'hDE)|(curr_ir == 8'hDB)|(curr_ir == 8'h83)|(curr_ir == 8'hD6)|(curr_ir == 8'h4E)|(curr_ir == 8'h7E)|(curr_ir == 8'hF6)|(curr_ir == 8'h21)|(curr_ir == 8'h61)|(curr_ir == 8'h71)|(curr_ir == 8'hB1)|(curr_ir == 8'h01)|(curr_ir == 8'hEE)|(curr_ir == 8'hFE)|(curr_ir == 8'h51)|(curr_ir == 8'h40)|(curr_ir == 8'h2F)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'h00)|(curr_ir == 8'h73)|(curr_ir == 8'h57)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hF3)|(curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'hE3)|(curr_ir == 8'h33)|(curr_ir == 8'h03)|(curr_ir == 8'h23)|(curr_ir == 8'h43)|(curr_ir == 8'hD3)|(curr_ir == 8'h73)|(curr_ir == 8'h13)|(curr_ir == 8'hC3)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hD3)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'hDE)|(curr_ir == 8'h1B)|(curr_ir == 8'hFE)|(curr_ir == 8'h73)|(curr_ir == 8'hFF)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'h1E)|(curr_ir == 8'h63)|(curr_ir == 8'hDF)|(curr_ir == 8'h7E)|(curr_ir == 8'hC3)|(curr_ir == 8'h5B)|(curr_ir == 8'h3E)|(curr_ir == 8'h00)|(curr_ir == 8'hE3)|(curr_ir == 8'hF3)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'hFB)|(curr_ir == 8'h1F)|(curr_ir == 8'h03)|(curr_ir == 8'hDB)|(curr_ir == 8'h53)|(curr_ir == 8'h5E)|(curr_ir == 8'h33)))|
	    ((curr_cycle == 0)))
		next_cycle = curr_cycle + 1;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h28)|(curr_ir == 8'h00)|(curr_ir == 8'h40)|(curr_ir == 8'h60)|(curr_ir == 8'h20)|(curr_ir == 8'h68)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h20)|(curr_ir == 8'h68)|(curr_ir == 8'h00)|(curr_ir == 8'h40)|(curr_ir == 8'h60)|(curr_ir == 8'h28)|(curr_ir == 8'h08)|(curr_ir == 8'h48)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h20)|(curr_ir == 8'h00)|(curr_ir == 8'h40)|(curr_ir == 8'h60)))|
	    ((curr_cycle == 5)&(curr_ir == 8'h40)))
		G_addr = curr_sp;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h8C)|(curr_ir == 8'h27)|(curr_ir == 8'hC7)|(curr_ir == 8'h94)|(curr_ir == 8'hE6)|(curr_ir == 8'hC6)|(curr_ir == 8'h07)|(curr_ir == 8'h8D)|(curr_ir == 8'h67)|(curr_ir == 8'h96)|(curr_ir == 8'h00)|(curr_ir == 8'h66)|(curr_ir == 8'h97)|(curr_ir == 8'h26)|(curr_ir == 8'hE7)|(curr_ir == 8'h46)|(curr_ir == 8'h06)|(curr_ir == 8'h8F)|(curr_ir == 8'h95)|(curr_ir == 8'h20)|(curr_ir == 8'h47)|(curr_ir == 8'h8E)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hFE)|(curr_ir == 8'hFF)|(curr_ir == 8'hDE)|(curr_ir == 8'hF3)|(curr_ir == 8'hDF)|(curr_ir == 8'hC3)|(curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'h23)|(curr_ir == 8'h5E)|(curr_ir == 8'hE3)|(curr_ir == 8'h33)|(curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'hFB)|(curr_ir == 8'h03)|(curr_ir == 8'h73)|(curr_ir == 8'hDB)|(curr_ir == 8'h43)|(curr_ir == 8'h13)|(curr_ir == 8'h1E)|(curr_ir == 8'hD3)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hE7)|(curr_ir == 8'h46)|(curr_ir == 8'hD7)|(curr_ir == 8'h37)|(curr_ir == 8'hD6)|(curr_ir == 8'h4E)|(curr_ir == 8'hF6)|(curr_ir == 8'hC6)|(curr_ir == 8'h9D)|(curr_ir == 8'h17)|(curr_ir == 8'h4F)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'h0E)|(curr_ir == 8'hCF)|(curr_ir == 8'h20)|(curr_ir == 8'hEE)|(curr_ir == 8'h16)|(curr_ir == 8'h77)|(curr_ir == 8'hCE)|(curr_ir == 8'hF7)|(curr_ir == 8'h26)|(curr_ir == 8'h99)|(curr_ir == 8'h66)|(curr_ir == 8'hC7)|(curr_ir == 8'h2E)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'h6F)|(curr_ir == 8'h2F)|(curr_ir == 8'h06)|(curr_ir == 8'h00)|(curr_ir == 8'hEF)|(curr_ir == 8'h0F)|(curr_ir == 8'h56)|(curr_ir == 8'h57)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h3E)|(curr_ir == 8'h0E)|(curr_ir == 8'hDB)|(curr_ir == 8'h6E)|(curr_ir == 8'hCF)|(curr_ir == 8'h1F)|(curr_ir == 8'h83)|(curr_ir == 8'h5E)|(curr_ir == 8'hEF)|(curr_ir == 8'h2E)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h91)|(curr_ir == 8'hFF)|(curr_ir == 8'hDE)|(curr_ir == 8'h4E)|(curr_ir == 8'h1B)|(curr_ir == 8'h1E)|(curr_ir == 8'h56)|(curr_ir == 8'hDF)|(curr_ir == 8'hF6)|(curr_ir == 8'h81)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'hF7)|(curr_ir == 8'hD6)|(curr_ir == 8'hD7)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h7E)|(curr_ir == 8'h16)|(curr_ir == 8'h5B)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'hFB)|(curr_ir == 8'hCE)))|
	    ((curr_cycle == 7)&((curr_ir == 8'hE3)|(curr_ir == 8'hD3)|(curr_ir == 8'hF3)|(curr_ir == 8'hC3)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h87)|(curr_ir == 8'h00)|(curr_ir == 8'h85)|(curr_ir == 8'h86)|(curr_ir == 8'h84)|(curr_ir == 8'h08)|(curr_ir == 8'h48)))|
	    ((curr_cycle == 1)&(curr_ir == 8'hCB)))
		G_rdwr = 0;
	
	if (((curr_cycle == 2)&(curr_ir == 8'h00))|
	    ((curr_cycle == 3)&(curr_ir == 8'h20)))
		G_wr_data = curr_pch;
	
	if (((curr_cycle == 2)&((curr_ir == 8'h00)|(curr_ir == 8'h08)|(curr_ir == 8'h48)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h00)|(curr_ir == 8'h20)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h20)|(curr_ir == 8'h00))))
		next_s = curr_s - 1;
	
	if (((curr_cycle == 3)&(curr_ir == 8'h00))|
	    ((curr_cycle == 4)&(curr_ir == 8'h20)))
		G_wr_data = curr_pcl;
	
	if (((curr_cycle == 4)&(curr_ir == 8'h00)))
		G_wr_data = curr_p | (is_soft_brk ? B_mask : 8'h00);
	
	if (((curr_cycle == 4)&(curr_ir == 8'h00)))
		next_p[I_bit] = irq_p | curr_p[I_bit];
	
	if (((curr_cycle == 5)&(curr_ir == 8'h00)))
		G_addr = vec_addr_lo;
	
	if (((curr_cycle == 1)&((curr_ir == 8'hD1)|(curr_ir == 8'hD7)|(curr_ir == 8'hC7)|(curr_ir == 8'hF5)|(curr_ir == 8'h34)|(curr_ir == 8'h95)|(curr_ir == 8'h85)|(curr_ir == 8'hC5)|(curr_ir == 8'h86)|(curr_ir == 8'h14)|(curr_ir == 8'h65)|(curr_ir == 8'hC6)|(curr_ir == 8'h17)|(curr_ir == 8'h11)|(curr_ir == 8'h53)|(curr_ir == 8'hB4)|(curr_ir == 8'hCD)|(curr_ir == 8'h20)|(curr_ir == 8'hEE)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h8E)|(curr_ir == 8'h84)|(curr_ir == 8'hCE)|(curr_ir == 8'h0F)|(curr_ir == 8'h2C)|(curr_ir == 8'h35)|(curr_ir == 8'hED)|(curr_ir == 8'h2E)|(curr_ir == 8'h66)|(curr_ir == 8'h54)|(curr_ir == 8'h73)|(curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'h57)|(curr_ir == 8'h94)|(curr_ir == 8'h25)|(curr_ir == 8'h6E)|(curr_ir == 8'hCF)|(curr_ir == 8'hE6)|(curr_ir == 8'h2D)|(curr_ir == 8'h55)|(curr_ir == 8'hB6)|(curr_ir == 8'h8D)|(curr_ir == 8'h07)|(curr_ir == 8'hAC)|(curr_ir == 8'h2F)|(curr_ir == 8'h06)|(curr_ir == 8'hE4)|(curr_ir == 8'hF1)|(curr_ir == 8'hD5)|(curr_ir == 8'h26)|(curr_ir == 8'h37)|(curr_ir == 8'h4E)|(curr_ir == 8'h05)|(curr_ir == 8'hA5)|(curr_ir == 8'hEF)|(curr_ir == 8'hD3)|(curr_ir == 8'h24)|(curr_ir == 8'h6D)|(curr_ir == 8'h31)|(curr_ir == 8'h4C)|(curr_ir == 8'hB7)|(curr_ir == 8'hC4)|(curr_ir == 8'h15)|(curr_ir == 8'h91)|(curr_ir == 8'h97)|(curr_ir == 8'h87)|(curr_ir == 8'h75)|(curr_ir == 8'hB5)|(curr_ir == 8'hCC)|(curr_ir == 8'h13)|(curr_ir == 8'hA6)|(curr_ir == 8'hD4)|(curr_ir == 8'h76)|(curr_ir == 8'h4D)|(curr_ir == 8'h74)|(curr_ir == 8'h64)|(curr_ir == 8'h71)|(curr_ir == 8'hAE)|(curr_ir == 8'hA4)|(curr_ir == 8'h0C)|(curr_ir == 8'h27)|(curr_ir == 8'hB1)|(curr_ir == 8'hAF)|(curr_ir == 8'h44)|(curr_ir == 8'hF6)|(curr_ir == 8'h47)|(curr_ir == 8'hEC)|(curr_ir == 8'h56)|(curr_ir == 8'h6F)|(curr_ir == 8'hA7)|(curr_ir == 8'hAD)|(curr_ir == 8'hE7)|(curr_ir == 8'h16)|(curr_ir == 8'hF4)|(curr_ir == 8'h46)|(curr_ir == 8'hE5)|(curr_ir == 8'h36)|(curr_ir == 8'h51)|(curr_ir == 8'h0D)|(curr_ir == 8'h4F)|(curr_ir == 8'h45)|(curr_ir == 8'h8F)|(curr_ir == 8'h96)|(curr_ir == 8'hF7)|(curr_ir == 8'h8C)|(curr_ir == 8'hB3)|(curr_ir == 8'h04)|(curr_ir == 8'hD6)|(curr_ir == 8'hF3)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h01)|(curr_ir == 8'h23)|(curr_ir == 8'hA3)|(curr_ir == 8'hE3)|(curr_ir == 8'hA1)|(curr_ir == 8'h83)|(curr_ir == 8'h41)|(curr_ir == 8'h63)|(curr_ir == 8'h6C)|(curr_ir == 8'h43)|(curr_ir == 8'h61)|(curr_ir == 8'hE1)|(curr_ir == 8'hC3)|(curr_ir == 8'h21)|(curr_ir == 8'h81)|(curr_ir == 8'hC1)|(curr_ir == 8'h03)))|
	    ((curr_cycle == 5)&(curr_ir == 8'h00)))
		next_adl = G_rd_data;
	
	if (((curr_cycle == 6)&(curr_ir == 8'h00)))
		G_addr = vec_addr_hi;
	
	if (((curr_cycle == 2)&((curr_ir == 8'hCD)|(curr_ir == 8'hCF)|(curr_ir == 8'h8E)|(curr_ir == 8'h4F)|(curr_ir == 8'h2D)|(curr_ir == 8'h8F)|(curr_ir == 8'hCC)|(curr_ir == 8'h8D)|(curr_ir == 8'hAC)|(curr_ir == 8'h2F)|(curr_ir == 8'hEE)|(curr_ir == 8'hCE)|(curr_ir == 8'h0D)|(curr_ir == 8'h8C)|(curr_ir == 8'h4D)|(curr_ir == 8'hAF)|(curr_ir == 8'h4E)|(curr_ir == 8'h2C)|(curr_ir == 8'h0F)|(curr_ir == 8'hAE)|(curr_ir == 8'hEF)|(curr_ir == 8'hED)|(curr_ir == 8'h2E)|(curr_ir == 8'h0C)|(curr_ir == 8'h6D)|(curr_ir == 8'hAD)|(curr_ir == 8'h6E)|(curr_ir == 8'h4C)|(curr_ir == 8'h6F)|(curr_ir == 8'h0E)|(curr_ir == 8'hEC)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h6C)|(curr_ir == 8'h43)|(curr_ir == 8'h21)|(curr_ir == 8'h81)|(curr_ir == 8'h61)|(curr_ir == 8'hC1)|(curr_ir == 8'h23)|(curr_ir == 8'h83)|(curr_ir == 8'h41)|(curr_ir == 8'hA3)|(curr_ir == 8'h03)|(curr_ir == 8'hE1)|(curr_ir == 8'hE3)|(curr_ir == 8'hA1)|(curr_ir == 8'h01)|(curr_ir == 8'h63)|(curr_ir == 8'hC3)))|
	    ((curr_cycle == 5)&(curr_ir == 8'h20))|
	    ((curr_cycle == 6)&(curr_ir == 8'h00)))
		next_adh = G_rd_data;
	
	if (((curr_cycle == 5)&(curr_ir == 8'h20))|
	    ((curr_cycle == 6)&(curr_ir == 8'h00))|
	    ((curr_cycle == 2)&(curr_ir == 8'h4C))|
	    ((curr_cycle == 4)&(curr_ir == 8'h6C)))
		{next_pch, next_pcl} = next_ad;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h0F)|(curr_ir == 8'h57)|(curr_ir == 8'h01)|(curr_ir == 8'h0E)|(curr_ir == 8'hA1)|(curr_ir == 8'h6E)|(curr_ir == 8'hCF)|(curr_ir == 8'h83)|(curr_ir == 8'hF1)|(curr_ir == 8'h60)|(curr_ir == 8'h40)|(curr_ir == 8'hEF)|(curr_ir == 8'h2E)|(curr_ir == 8'h31)|(curr_ir == 8'h91)|(curr_ir == 8'h2F)|(curr_ir == 8'h41)|(curr_ir == 8'h4E)|(curr_ir == 8'hE1)|(curr_ir == 8'h56)|(curr_ir == 8'hF6)|(curr_ir == 8'h81)|(curr_ir == 8'hC1)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'h71)|(curr_ir == 8'hF7)|(curr_ir == 8'h37)|(curr_ir == 8'hD6)|(curr_ir == 8'hD1)|(curr_ir == 8'hD7)|(curr_ir == 8'h6F)|(curr_ir == 8'hB1)|(curr_ir == 8'h20)|(curr_ir == 8'h16)|(curr_ir == 8'h21)|(curr_ir == 8'h11)|(curr_ir == 8'h17)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h4F)|(curr_ir == 8'hEE)|(curr_ir == 8'h77)|(curr_ir == 8'hB3)|(curr_ir == 8'hCE)|(curr_ir == 8'hA3)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h8C)|(curr_ir == 8'hED)|(curr_ir == 8'h70)|(curr_ir == 8'h34)|(curr_ir == 8'h94)|(curr_ir == 8'h50)|(curr_ir == 8'hF5)|(curr_ir == 8'hB6)|(curr_ir == 8'h8D)|(curr_ir == 8'hF4)|(curr_ir == 8'h35)|(curr_ir == 8'h10)|(curr_ir == 8'h96)|(curr_ir == 8'hAF)|(curr_ir == 8'h97)|(curr_ir == 8'h75)|(curr_ir == 8'h2D)|(curr_ir == 8'hCC)|(curr_ir == 8'hB0)|(curr_ir == 8'hCD)|(curr_ir == 8'h68)|(curr_ir == 8'hAC)|(curr_ir == 8'h90)|(curr_ir == 8'h74)|(curr_ir == 8'h28)|(curr_ir == 8'hAE)|(curr_ir == 8'hD5)|(curr_ir == 8'hB7)|(curr_ir == 8'hAD)|(curr_ir == 8'h15)|(curr_ir == 8'hB4)|(curr_ir == 8'h55)|(curr_ir == 8'hB5)|(curr_ir == 8'h8F)|(curr_ir == 8'hF0)|(curr_ir == 8'hD4)|(curr_ir == 8'h4D)|(curr_ir == 8'h0C)|(curr_ir == 8'h6D)|(curr_ir == 8'h95)|(curr_ir == 8'h30)|(curr_ir == 8'hEC)|(curr_ir == 8'h14)|(curr_ir == 8'hD0)|(curr_ir == 8'h8E)|(curr_ir == 8'h0D)|(curr_ir == 8'h2C)|(curr_ir == 8'h54)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h18)|(curr_ir == 8'h5A)|(curr_ir == 8'h88)|(curr_ir == 8'hC0)|(curr_ir == 8'h49)|(curr_ir == 8'hA0)|(curr_ir == 8'hA2)|(curr_ir == 8'hC9)|(curr_ir == 8'hFA)|(curr_ir == 8'h4A)|(curr_ir == 8'hAB)|(curr_ir == 8'hB8)|(curr_ir == 8'h09)|(curr_ir == 8'hEB)|(curr_ir == 8'h1A)|(curr_ir == 8'hF8)|(curr_ir == 8'h69)|(curr_ir == 8'hA9)|(curr_ir == 8'h9A)|(curr_ir == 8'hCA)|(curr_ir == 8'hDA)|(curr_ir == 8'h38)|(curr_ir == 8'hC8)|(curr_ir == 8'h6A)|(curr_ir == 8'hCB)|(curr_ir == 8'h58)|(curr_ir == 8'h98)|(curr_ir == 8'h89)|(curr_ir == 8'hEA)|(curr_ir == 8'hE0)|(curr_ir == 8'h3A)|(curr_ir == 8'h7A)|(curr_ir == 8'hC2)|(curr_ir == 8'h2A)|(curr_ir == 8'h80)|(curr_ir == 8'hE9)|(curr_ir == 8'hBA)|(curr_ir == 8'h0A)|(curr_ir == 8'hAA)|(curr_ir == 8'hE2)|(curr_ir == 8'hD8)|(curr_ir == 8'hE8)|(curr_ir == 8'h29)|(curr_ir == 8'h78)|(curr_ir == 8'hA8)|(curr_ir == 8'h8A)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hFE)|(curr_ir == 8'hFF)|(curr_ir == 8'hDE)|(curr_ir == 8'h1F)|(curr_ir == 8'h3F)|(curr_ir == 8'hDF)|(curr_ir == 8'h5E)|(curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'hFB)|(curr_ir == 8'h5B)|(curr_ir == 8'h00)|(curr_ir == 8'h1B)|(curr_ir == 8'h3B)|(curr_ir == 8'hDB)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h1E)|(curr_ir == 8'h7F)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hE7)|(curr_ir == 8'hD9)|(curr_ir == 8'h39)|(curr_ir == 8'h46)|(curr_ir == 8'hFD)|(curr_ir == 8'hBE)|(curr_ir == 8'h27)|(curr_ir == 8'hF9)|(curr_ir == 8'hB9)|(curr_ir == 8'hC6)|(curr_ir == 8'h9D)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'h5C)|(curr_ir == 8'hFC)|(curr_ir == 8'h19)|(curr_ir == 8'h79)|(curr_ir == 8'hDC)|(curr_ir == 8'h3C)|(curr_ir == 8'h07)|(curr_ir == 8'hBC)|(curr_ir == 8'hBF)|(curr_ir == 8'h26)|(curr_ir == 8'h99)|(curr_ir == 8'h66)|(curr_ir == 8'h7D)|(curr_ir == 8'hC7)|(curr_ir == 8'hBD)|(curr_ir == 8'hE6)|(curr_ir == 8'h6C)|(curr_ir == 8'h06)|(curr_ir == 8'h1D)|(curr_ir == 8'h5D)|(curr_ir == 8'h67)|(curr_ir == 8'h7C)|(curr_ir == 8'h1C)|(curr_ir == 8'hDD)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h33)|(curr_ir == 8'hE3)|(curr_ir == 8'hD3)|(curr_ir == 8'h73)|(curr_ir == 8'h63)|(curr_ir == 8'h43)|(curr_ir == 8'h13)|(curr_ir == 8'hF3)|(curr_ir == 8'hC3)|(curr_ir == 8'h03)|(curr_ir == 8'h53)|(curr_ir == 8'h23)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h04)|(curr_ir == 8'h44)|(curr_ir == 8'hA5)|(curr_ir == 8'h4C)|(curr_ir == 8'hC4)|(curr_ir == 8'h87)|(curr_ir == 8'h45)|(curr_ir == 8'hA6)|(curr_ir == 8'h64)|(curr_ir == 8'hA4)|(curr_ir == 8'h25)|(curr_ir == 8'h65)|(curr_ir == 8'hA7)|(curr_ir == 8'hC5)|(curr_ir == 8'h48)|(curr_ir == 8'hE5)|(curr_ir == 8'hE4)|(curr_ir == 8'h05)|(curr_ir == 8'h85)|(curr_ir == 8'h86)|(curr_ir == 8'h84)|(curr_ir == 8'h24)|(curr_ir == 8'h08))))
		next_cycle = 0;
	
	if (((curr_cycle == 1)&((curr_ir == 8'hD1)|(curr_ir == 8'h22)|(curr_ir == 8'hC7)|(curr_ir == 8'hD7)|(curr_ir == 8'h3F)|(curr_ir == 8'h50)|(curr_ir == 8'h3E)|(curr_ir == 8'h34)|(curr_ir == 8'hF5)|(curr_ir == 8'h7E)|(curr_ir == 8'h95)|(curr_ir == 8'h85)|(curr_ir == 8'h01)|(curr_ir == 8'h79)|(curr_ir == 8'hC5)|(curr_ir == 8'h3D)|(curr_ir == 8'h86)|(curr_ir == 8'h14)|(curr_ir == 8'hC3)|(curr_ir == 8'hD0)|(curr_ir == 8'h65)|(curr_ir == 8'h21)|(curr_ir == 8'h3C)|(curr_ir == 8'h11)|(curr_ir == 8'h17)|(curr_ir == 8'hC0)|(curr_ir == 8'h53)|(curr_ir == 8'hB4)|(curr_ir == 8'h49)|(curr_ir == 8'hC6)|(curr_ir == 8'h20)|(curr_ir == 8'hCD)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'hA0)|(curr_ir == 8'hFB)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h8E)|(curr_ir == 8'h84)|(curr_ir == 8'h5B)|(curr_ir == 8'hCE)|(curr_ir == 8'h1F)|(curr_ir == 8'h0F)|(curr_ir == 8'h2C)|(curr_ir == 8'h03)|(curr_ir == 8'hA2)|(curr_ir == 8'hB2)|(curr_ir == 8'hC9)|(curr_ir == 8'hBF)|(curr_ir == 8'h35)|(curr_ir == 8'h10)|(curr_ir == 8'hA3)|(curr_ir == 8'hF9)|(curr_ir == 8'hED)|(curr_ir == 8'hDD)|(curr_ir == 8'h2E)|(curr_ir == 8'h70)|(curr_ir == 8'h66)|(curr_ir == 8'h7D)|(curr_ir == 8'h54)|(curr_ir == 8'h73)|(curr_ir == 8'hBD)|(curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'h57)|(curr_ir == 8'h94)|(curr_ir == 8'h25)|(curr_ir == 8'hAB)|(curr_ir == 8'hA1)|(curr_ir == 8'h09)|(curr_ir == 8'hEB)|(curr_ir == 8'hDB)|(curr_ir == 8'h6E)|(curr_ir == 8'h92)|(curr_ir == 8'hCF)|(curr_ir == 8'hE6)|(curr_ir == 8'h7B)|(curr_ir == 8'hDC)|(curr_ir == 8'h2D)|(curr_ir == 8'h69)|(curr_ir == 8'h5F)|(curr_ir == 8'h55)|(curr_ir == 8'h6C)|(curr_ir == 8'hA9)|(curr_ir == 8'h43)|(curr_ir == 8'hB6)|(curr_ir == 8'h07)|(curr_ir == 8'h8D)|(curr_ir == 8'h83)|(curr_ir == 8'hAC)|(curr_ir == 8'h2F)|(curr_ir == 8'h90)|(curr_ir == 8'h06)|(curr_ir == 8'hE4)|(curr_ir == 8'hF1)|(curr_ir == 8'h42)|(curr_ir == 8'h5D)|(curr_ir == 8'hBE)|(curr_ir == 8'hD5)|(curr_ir == 8'h26)|(curr_ir == 8'h41)|(curr_ir == 8'h1C)|(curr_ir == 8'h37)|(curr_ir == 8'hCB)|(curr_ir == 8'h5E)|(curr_ir == 8'h05)|(curr_ir == 8'h4E)|(curr_ir == 8'h12)|(curr_ir == 8'hA5)|(curr_ir == 8'h7C)|(curr_ir == 8'h99)|(curr_ir == 8'hEF)|(curr_ir == 8'h89)|(curr_ir == 8'hD3)|(curr_ir == 8'h24)|(curr_ir == 8'h6D)|(curr_ir == 8'h3B)|(curr_ir == 8'hE0)|(curr_ir == 8'h31)|(curr_ir == 8'h4C)|(curr_ir == 8'hB7)|(curr_ir == 8'hC4)|(curr_ir == 8'h59)|(curr_ir == 8'h15)|(curr_ir == 8'h30)|(curr_ir == 8'h91)|(curr_ir == 8'h97)|(curr_ir == 8'h87)|(curr_ir == 8'hF2)|(curr_ir == 8'h75)|(curr_ir == 8'hFF)|(curr_ir == 8'h82)|(curr_ir == 8'hDE)|(curr_ir == 8'hB5)|(curr_ir == 8'hCC)|(curr_ir == 8'hD2)|(curr_ir == 8'h1D)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'hC2)|(curr_ir == 8'hD9)|(curr_ir == 8'hB0)|(curr_ir == 8'hA6)|(curr_ir == 8'h39)|(curr_ir == 8'hF0)|(curr_ir == 8'hFD)|(curr_ir == 8'hD4)|(curr_ir == 8'h76)|(curr_ir == 8'h32)|(curr_ir == 8'h4D)|(curr_ir == 8'h80)|(curr_ir == 8'hE1)|(curr_ir == 8'h74)|(curr_ir == 8'h64)|(curr_ir == 8'h71)|(curr_ir == 8'h1E)|(curr_ir == 8'hA4)|(curr_ir == 8'hAE)|(curr_ir == 8'h0C)|(curr_ir == 8'h27)|(curr_ir == 8'h02)|(curr_ir == 8'hB1)|(curr_ir == 8'hAF)|(curr_ir == 8'h44)|(curr_ir == 8'h19)|(curr_ir == 8'h1B)|(curr_ir == 8'hE9)|(curr_ir == 8'hDF)|(curr_ir == 8'hF6)|(curr_ir == 8'h72)|(curr_ir == 8'h47)|(curr_ir == 8'h62)|(curr_ir == 8'hEC)|(curr_ir == 8'h7F)|(curr_ir == 8'h56)|(curr_ir == 8'h6F)|(curr_ir == 8'h63)|(curr_ir == 8'hB9)|(curr_ir == 8'hA7)|(curr_ir == 8'hAD)|(curr_ir == 8'h9D)|(curr_ir == 8'hE3)|(curr_ir == 8'hE7)|(curr_ir == 8'h81)|(curr_ir == 8'h16)|(curr_ir == 8'hF4)|(curr_ir == 8'hC1)|(curr_ir == 8'hE2)|(curr_ir == 8'h29)|(curr_ir == 8'h46)|(curr_ir == 8'h61)|(curr_ir == 8'h36)|(curr_ir == 8'h51)|(curr_ir == 8'h0D)|(curr_ir == 8'hBC)|(curr_ir == 8'hE5)|(curr_ir == 8'h4F)|(curr_ir == 8'h45)|(curr_ir == 8'hFC)|(curr_ir == 8'h5C)|(curr_ir == 8'h52)|(curr_ir == 8'h8F)|(curr_ir == 8'h96)|(curr_ir == 8'hF7)|(curr_ir == 8'h8C)|(curr_ir == 8'hB3)|(curr_ir == 8'h04)|(curr_ir == 8'hD6)|(curr_ir == 8'hF3)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h5F)|(curr_ir == 8'h6C)|(curr_ir == 8'h8F)|(curr_ir == 8'h8D)|(curr_ir == 8'hAC)|(curr_ir == 8'h2F)|(curr_ir == 8'h1D)|(curr_ir == 8'h5D)|(curr_ir == 8'h4E)|(curr_ir == 8'h3F)|(curr_ir == 8'h7C)|(curr_ir == 8'h1E)|(curr_ir == 8'h7F)|(curr_ir == 8'h0C)|(curr_ir == 8'h6D)|(curr_ir == 8'h59)|(curr_ir == 8'hDF)|(curr_ir == 8'h3D)|(curr_ir == 8'hEC)|(curr_ir == 8'hFF)|(curr_ir == 8'hFE)|(curr_ir == 8'h4F)|(curr_ir == 8'hCC)|(curr_ir == 8'h5C)|(curr_ir == 8'hD9)|(curr_ir == 8'hCE)|(curr_ir == 8'hDE)|(curr_ir == 8'h1F)|(curr_ir == 8'h0D)|(curr_ir == 8'hFC)|(curr_ir == 8'h4D)|(curr_ir == 8'hAE)|(curr_ir == 8'h19)|(curr_ir == 8'h6F)|(curr_ir == 8'hB9)|(curr_ir == 8'h9D)|(curr_ir == 8'h8E)|(curr_ir == 8'hBC)|(curr_ir == 8'h5E)|(curr_ir == 8'hEE)|(curr_ir == 8'h8C)|(curr_ir == 8'h99)|(curr_ir == 8'h2C)|(curr_ir == 8'hEF)|(curr_ir == 8'hED)|(curr_ir == 8'h3E)|(curr_ir == 8'h2E)|(curr_ir == 8'hDD)|(curr_ir == 8'h3B)|(curr_ir == 8'h7E)|(curr_ir == 8'h6E)|(curr_ir == 8'h7B)|(curr_ir == 8'h79)|(curr_ir == 8'h0E)|(curr_ir == 8'h3C)|(curr_ir == 8'hDB)|(curr_ir == 8'hCD)|(curr_ir == 8'hCF)|(curr_ir == 8'h39)|(curr_ir == 8'h2D)|(curr_ir == 8'hFD)|(curr_ir == 8'hFB)|(curr_ir == 8'h5B)|(curr_ir == 8'hBE)|(curr_ir == 8'hAF)|(curr_ir == 8'hBF)|(curr_ir == 8'h1B)|(curr_ir == 8'h0F)|(curr_ir == 8'h1C)|(curr_ir == 8'h7D)|(curr_ir == 8'hF9)|(curr_ir == 8'hBD)|(curr_ir == 8'hAD)|(curr_ir == 8'hDC)))|
	    ((curr_cycle == 5)&(curr_ir == 8'h60)))
		{next_pch, next_pcl} = curr_pc + 1;
	
	if (((curr_cycle == 1)&((curr_ir == 8'hA1)|(curr_ir == 8'h01)|(curr_ir == 8'hC1)|(curr_ir == 8'h43)|(curr_ir == 8'h03)|(curr_ir == 8'h63)|(curr_ir == 8'h23)|(curr_ir == 8'hE1)|(curr_ir == 8'h41)|(curr_ir == 8'h83)|(curr_ir == 8'hC3)|(curr_ir == 8'h61)|(curr_ir == 8'hA3)|(curr_ir == 8'h21)|(curr_ir == 8'hE3)|(curr_ir == 8'h81))))
		next_bah = 0;
	
	if (((curr_cycle == 1)&((curr_ir == 8'hDD)|(curr_ir == 8'h7C)|(curr_ir == 8'h3F)|(curr_ir == 8'h19)|(curr_ir == 8'h1B)|(curr_ir == 8'h7D)|(curr_ir == 8'h99)|(curr_ir == 8'hF9)|(curr_ir == 8'h3E)|(curr_ir == 8'hDF)|(curr_ir == 8'hBD)|(curr_ir == 8'h7E)|(curr_ir == 8'h3B)|(curr_ir == 8'hA1)|(curr_ir == 8'h7F)|(curr_ir == 8'h01)|(curr_ir == 8'h59)|(curr_ir == 8'h79)|(curr_ir == 8'hDB)|(curr_ir == 8'h63)|(curr_ir == 8'hB9)|(curr_ir == 8'h3D)|(curr_ir == 8'hC3)|(curr_ir == 8'h9D)|(curr_ir == 8'h7B)|(curr_ir == 8'hDC)|(curr_ir == 8'h21)|(curr_ir == 8'h3C)|(curr_ir == 8'hFF)|(curr_ir == 8'h81)|(curr_ir == 8'h5F)|(curr_ir == 8'hDE)|(curr_ir == 8'h6C)|(curr_ir == 8'hC1)|(curr_ir == 8'h43)|(curr_ir == 8'hFE)|(curr_ir == 8'h1D)|(curr_ir == 8'h23)|(curr_ir == 8'hFB)|(curr_ir == 8'h83)|(curr_ir == 8'hD9)|(curr_ir == 8'h61)|(curr_ir == 8'hBC)|(curr_ir == 8'h5B)|(curr_ir == 8'h39)|(curr_ir == 8'hFC)|(curr_ir == 8'h1F)|(curr_ir == 8'h5C)|(curr_ir == 8'hFD)|(curr_ir == 8'h5D)|(curr_ir == 8'hBE)|(curr_ir == 8'h03)|(curr_ir == 8'hE1)|(curr_ir == 8'hBF)|(curr_ir == 8'h41)|(curr_ir == 8'h1C)|(curr_ir == 8'h5E)|(curr_ir == 8'hA3)|(curr_ir == 8'hE3)|(curr_ir == 8'h1E)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h11)|(curr_ir == 8'h51)|(curr_ir == 8'hB3)|(curr_ir == 8'h13)|(curr_ir == 8'hF1)|(curr_ir == 8'hF3)|(curr_ir == 8'h71)|(curr_ir == 8'hD1)|(curr_ir == 8'h33)|(curr_ir == 8'hB1)|(curr_ir == 8'h73)|(curr_ir == 8'h91)|(curr_ir == 8'hD3)|(curr_ir == 8'h31)|(curr_ir == 8'h53))))
		next_bal = G_rd_data;
	
	if (((curr_cycle == 2)&((curr_ir == 8'h81)|(curr_ir == 8'h23)|(curr_ir == 8'h43)|(curr_ir == 8'h83)|(curr_ir == 8'h61)|(curr_ir == 8'hC1)|(curr_ir == 8'hE1)|(curr_ir == 8'h41)|(curr_ir == 8'hA3)|(curr_ir == 8'h03)|(curr_ir == 8'hE3)|(curr_ir == 8'hC3)|(curr_ir == 8'hA1)|(curr_ir == 8'h01)|(curr_ir == 8'h63)|(curr_ir == 8'h21)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hE1)|(curr_ir == 8'h41)|(curr_ir == 8'hA3)|(curr_ir == 8'h01)|(curr_ir == 8'h63)|(curr_ir == 8'hE3)|(curr_ir == 8'hC3)|(curr_ir == 8'hA1)|(curr_ir == 8'h21)|(curr_ir == 8'h23)|(curr_ir == 8'h6C)|(curr_ir == 8'h43)|(curr_ir == 8'h81)|(curr_ir == 8'h61)|(curr_ir == 8'hC1)|(curr_ir == 8'h83)|(curr_ir == 8'h03)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h6C)|(curr_ir == 8'h43)|(curr_ir == 8'h21)|(curr_ir == 8'h81)|(curr_ir == 8'h61)|(curr_ir == 8'hC1)|(curr_ir == 8'h23)|(curr_ir == 8'h83)|(curr_ir == 8'h41)|(curr_ir == 8'hA3)|(curr_ir == 8'h03)|(curr_ir == 8'hE1)|(curr_ir == 8'hE3)|(curr_ir == 8'hA1)|(curr_ir == 8'h01)|(curr_ir == 8'h63)|(curr_ir == 8'hC3))))
		G_addr = curr_ba;
	
	if (((curr_cycle == 2)&((curr_ir == 8'h81)|(curr_ir == 8'hA1)|(curr_ir == 8'h01)|(curr_ir == 8'h23)|(curr_ir == 8'hA3)|(curr_ir == 8'hC3)|(curr_ir == 8'h43)|(curr_ir == 8'h63)|(curr_ir == 8'hE1)|(curr_ir == 8'h41)|(curr_ir == 8'h83)|(curr_ir == 8'hE3)|(curr_ir == 8'h61)|(curr_ir == 8'hC1)|(curr_ir == 8'h21)|(curr_ir == 8'h03))))
		next_bal = curr_bal + curr_x;
	
	if (((curr_cycle == 3)&((curr_ir == 8'hE1)|(curr_ir == 8'h63)|(curr_ir == 8'h41)|(curr_ir == 8'h83)|(curr_ir == 8'h23)|(curr_ir == 8'h6C)|(curr_ir == 8'hA1)|(curr_ir == 8'h43)|(curr_ir == 8'h03)|(curr_ir == 8'hA3)|(curr_ir == 8'hE3)|(curr_ir == 8'h81)|(curr_ir == 8'hC3)|(curr_ir == 8'h01)|(curr_ir == 8'h61)|(curr_ir == 8'hC1)|(curr_ir == 8'h21))))
		next_bal = curr_bal + 1;
	
	if (((curr_cycle == 3)&((curr_ir == 8'hC7)|(curr_ir == 8'h33)|(curr_ir == 8'h0E)|(curr_ir == 8'h53)|(curr_ir == 8'hC6)|(curr_ir == 8'hB6)|(curr_ir == 8'h67)|(curr_ir == 8'h66)|(curr_ir == 8'h56)|(curr_ir == 8'hCD)|(curr_ir == 8'hAE)|(curr_ir == 8'h26)|(curr_ir == 8'h31)|(curr_ir == 8'hAD)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'h06)|(curr_ir == 8'h4D)|(curr_ir == 8'h6D)|(curr_ir == 8'hEC)|(curr_ir == 8'h0D)|(curr_ir == 8'h8C)|(curr_ir == 8'h34)|(curr_ir == 8'hD1)|(curr_ir == 8'h94)|(curr_ir == 8'hF5)|(curr_ir == 8'h6F)|(curr_ir == 8'h17)|(curr_ir == 8'h07)|(curr_ir == 8'hF4)|(curr_ir == 8'hAF)|(curr_ir == 8'hEF)|(curr_ir == 8'hD3)|(curr_ir == 8'h0F)|(curr_ir == 8'hB7)|(curr_ir == 8'hE7)|(curr_ir == 8'h4F)|(curr_ir == 8'h4E)|(curr_ir == 8'hB1)|(curr_ir == 8'h95)|(curr_ir == 8'hF6)|(curr_ir == 8'h51)|(curr_ir == 8'h2C)|(curr_ir == 8'h71)|(curr_ir == 8'hED)|(curr_ir == 8'hD6)|(curr_ir == 8'h11)|(curr_ir == 8'h8D)|(curr_ir == 8'hEE)|(curr_ir == 8'h35)|(curr_ir == 8'h97)|(curr_ir == 8'hCC)|(curr_ir == 8'h37)|(curr_ir == 8'h73)|(curr_ir == 8'h57)|(curr_ir == 8'h46)|(curr_ir == 8'h2F)|(curr_ir == 8'h13)|(curr_ir == 8'h8F)|(curr_ir == 8'hD4)|(curr_ir == 8'h76)|(curr_ir == 8'hCF)|(curr_ir == 8'h47)|(curr_ir == 8'h8E)|(curr_ir == 8'hCE)|(curr_ir == 8'h36)|(curr_ir == 8'hF7)|(curr_ir == 8'h27)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'h16)|(curr_ir == 8'hF1)|(curr_ir == 8'h96)|(curr_ir == 8'h2E)|(curr_ir == 8'h91)|(curr_ir == 8'h75)|(curr_ir == 8'h2D)|(curr_ir == 8'hAC)|(curr_ir == 8'h74)|(curr_ir == 8'hD5)|(curr_ir == 8'hB4)|(curr_ir == 8'hB5)|(curr_ir == 8'hB3)|(curr_ir == 8'hF3)|(curr_ir == 8'hD7)|(curr_ir == 8'h0C)|(curr_ir == 8'h14)|(curr_ir == 8'h77)|(curr_ir == 8'h54)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h57)|(curr_ir == 8'h83)|(curr_ir == 8'hEF)|(curr_ir == 8'hD3)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'hDE)|(curr_ir == 8'h4E)|(curr_ir == 8'h1B)|(curr_ir == 8'hF6)|(curr_ir == 8'h71)|(curr_ir == 8'hD6)|(curr_ir == 8'hB1)|(curr_ir == 8'h21)|(curr_ir == 8'h11)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'h01)|(curr_ir == 8'h73)|(curr_ir == 8'hFF)|(curr_ir == 8'h2F)|(curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'h1E)|(curr_ir == 8'h63)|(curr_ir == 8'hDF)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'hF7)|(curr_ir == 8'h37)|(curr_ir == 8'h7E)|(curr_ir == 8'h16)|(curr_ir == 8'hC3)|(curr_ir == 8'h5B)|(curr_ir == 8'h4F)|(curr_ir == 8'hCE)|(curr_ir == 8'h3E)|(curr_ir == 8'hA1)|(curr_ir == 8'h6E)|(curr_ir == 8'hF1)|(curr_ir == 8'h2E)|(curr_ir == 8'h91)|(curr_ir == 8'h41)|(curr_ir == 8'hF3)|(curr_ir == 8'hE3)|(curr_ir == 8'hD7)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h6F)|(curr_ir == 8'hFB)|(curr_ir == 8'h77)|(curr_ir == 8'hB3)|(curr_ir == 8'hA3)|(curr_ir == 8'h1F)|(curr_ir == 8'h0F)|(curr_ir == 8'h03)|(curr_ir == 8'h0E)|(curr_ir == 8'hDB)|(curr_ir == 8'h53)|(curr_ir == 8'hCF)|(curr_ir == 8'h5E)|(curr_ir == 8'h33)|(curr_ir == 8'h31)|(curr_ir == 8'hE1)|(curr_ir == 8'h56)|(curr_ir == 8'h81)|(curr_ir == 8'hC1)|(curr_ir == 8'hD1)|(curr_ir == 8'h17)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h46)|(curr_ir == 8'hD7)|(curr_ir == 8'h37)|(curr_ir == 8'h27)|(curr_ir == 8'hC6)|(curr_ir == 8'hFF)|(curr_ir == 8'h5B)|(curr_ir == 8'h4F)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'h3E)|(curr_ir == 8'hDF)|(curr_ir == 8'hCF)|(curr_ir == 8'h16)|(curr_ir == 8'hCE)|(curr_ir == 8'hF7)|(curr_ir == 8'h99)|(curr_ir == 8'h7D)|(curr_ir == 8'hBD)|(curr_ir == 8'h2E)|(curr_ir == 8'h6E)|(curr_ir == 8'hE6)|(curr_ir == 8'h1D)|(curr_ir == 8'h5D)|(curr_ir == 8'h1C)|(curr_ir == 8'hF9)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h1F)|(curr_ir == 8'hFC)|(curr_ir == 8'h1E)|(curr_ir == 8'h0E)|(curr_ir == 8'h77)|(curr_ir == 8'hBC)|(curr_ir == 8'h5E)|(curr_ir == 8'h26)|(curr_ir == 8'h66)|(curr_ir == 8'hC7)|(curr_ir == 8'h06)|(curr_ir == 8'hFB)|(curr_ir == 8'h67)|(curr_ir == 8'h56)|(curr_ir == 8'hD9)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'hBE)|(curr_ir == 8'hB9)|(curr_ir == 8'h9D)|(curr_ir == 8'h17)|(curr_ir == 8'h5C)|(curr_ir == 8'hDC)|(curr_ir == 8'h3C)|(curr_ir == 8'h07)|(curr_ir == 8'hBF)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h6F)|(curr_ir == 8'h5F)|(curr_ir == 8'h1B)|(curr_ir == 8'hEF)|(curr_ir == 8'h0F)|(curr_ir == 8'hDE)|(curr_ir == 8'hE7)|(curr_ir == 8'hDB)|(curr_ir == 8'hD6)|(curr_ir == 8'h4E)|(curr_ir == 8'h7E)|(curr_ir == 8'hF6)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'h19)|(curr_ir == 8'h79)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'h2F)|(curr_ir == 8'h7C)|(curr_ir == 8'hDD)|(curr_ir == 8'h57)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h1F)|(curr_ir == 8'hF3)|(curr_ir == 8'h3F)|(curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'h5E)|(curr_ir == 8'hE3)|(curr_ir == 8'h33)|(curr_ir == 8'hFB)|(curr_ir == 8'h5B)|(curr_ir == 8'h03)|(curr_ir == 8'hDB)|(curr_ir == 8'hFE)|(curr_ir == 8'h23)|(curr_ir == 8'h1B)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h43)|(curr_ir == 8'hD3)|(curr_ir == 8'hDE)|(curr_ir == 8'h73)|(curr_ir == 8'h13)|(curr_ir == 8'h1E)|(curr_ir == 8'hFF)|(curr_ir == 8'hDF)|(curr_ir == 8'hC3)|(curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'h7F)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hB7)|(curr_ir == 8'hE7)|(curr_ir == 8'hA6)|(curr_ir == 8'h71)|(curr_ir == 8'hD6)|(curr_ir == 8'hB1)|(curr_ir == 8'h95)|(curr_ir == 8'hF6)|(curr_ir == 8'hA7)|(curr_ir == 8'hC5)|(curr_ir == 8'h11)|(curr_ir == 8'hE5)|(curr_ir == 8'h51)|(curr_ir == 8'h35)|(curr_ir == 8'h96)|(curr_ir == 8'h85)|(curr_ir == 8'h84)|(curr_ir == 8'h74)|(curr_ir == 8'h73)|(curr_ir == 8'h57)|(curr_ir == 8'h24)|(curr_ir == 8'h46)|(curr_ir == 8'h13)|(curr_ir == 8'h37)|(curr_ir == 8'hD4)|(curr_ir == 8'h47)|(curr_ir == 8'h87)|(curr_ir == 8'h36)|(curr_ir == 8'h76)|(curr_ir == 8'hF7)|(curr_ir == 8'h27)|(curr_ir == 8'h25)|(curr_ir == 8'h65)|(curr_ir == 8'h16)|(curr_ir == 8'h05)|(curr_ir == 8'hE6)|(curr_ir == 8'hF1)|(curr_ir == 8'h91)|(curr_ir == 8'hB5)|(curr_ir == 8'hD5)|(curr_ir == 8'hF3)|(curr_ir == 8'hC4)|(curr_ir == 8'h14)|(curr_ir == 8'h75)|(curr_ir == 8'hB3)|(curr_ir == 8'h64)|(curr_ir == 8'hA4)|(curr_ir == 8'h53)|(curr_ir == 8'hD7)|(curr_ir == 8'hC7)|(curr_ir == 8'h33)|(curr_ir == 8'h86)|(curr_ir == 8'hC6)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h26)|(curr_ir == 8'h66)|(curr_ir == 8'h56)|(curr_ir == 8'h31)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'hB6)|(curr_ir == 8'h06)|(curr_ir == 8'h04)|(curr_ir == 8'h44)|(curr_ir == 8'hA5)|(curr_ir == 8'h45)|(curr_ir == 8'h34)|(curr_ir == 8'hF5)|(curr_ir == 8'h17)|(curr_ir == 8'hF4)|(curr_ir == 8'hE4)|(curr_ir == 8'hD1)|(curr_ir == 8'h97)|(curr_ir == 8'hB4)|(curr_ir == 8'h07)|(curr_ir == 8'h54)|(curr_ir == 8'h94)|(curr_ir == 8'hD3)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h73)|(curr_ir == 8'h63)|(curr_ir == 8'h13)|(curr_ir == 8'hC3)|(curr_ir == 8'hF3)|(curr_ir == 8'h03)|(curr_ir == 8'h53)|(curr_ir == 8'h33)|(curr_ir == 8'h23)|(curr_ir == 8'hD3)|(curr_ir == 8'hE3)|(curr_ir == 8'h43))))
		G_addr = curr_ad;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h0F)|(curr_ir == 8'h03)|(curr_ir == 8'h57)|(curr_ir == 8'h01)|(curr_ir == 8'h53)|(curr_ir == 8'hD3)|(curr_ir == 8'h31)|(curr_ir == 8'h43)|(curr_ir == 8'h2F)|(curr_ir == 8'h13)|(curr_ir == 8'h41)|(curr_ir == 8'hC1)|(curr_ir == 8'h37)|(curr_ir == 8'hD1)|(curr_ir == 8'hC3)|(curr_ir == 8'h21)|(curr_ir == 8'h11)|(curr_ir == 8'h17)|(curr_ir == 8'h51)|(curr_ir == 8'h4F)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hD6)|(curr_ir == 8'h0E)|(curr_ir == 8'h16)|(curr_ir == 8'h17)|(curr_ir == 8'hEE)|(curr_ir == 8'h35)|(curr_ir == 8'h56)|(curr_ir == 8'h2D)|(curr_ir == 8'hCC)|(curr_ir == 8'hCD)|(curr_ir == 8'h0F)|(curr_ir == 8'hD5)|(curr_ir == 8'h57)|(curr_ir == 8'h15)|(curr_ir == 8'h4F)|(curr_ir == 8'h55)|(curr_ir == 8'h4E)|(curr_ir == 8'hD7)|(curr_ir == 8'h4D)|(curr_ir == 8'hCF)|(curr_ir == 8'hF6)|(curr_ir == 8'hEC)|(curr_ir == 8'hCE)|(curr_ir == 8'h0D)|(curr_ir == 8'h2C)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hDE)|(curr_ir == 8'hD9)|(curr_ir == 8'hDB)|(curr_ir == 8'h39)|(curr_ir == 8'h27)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'h5B)|(curr_ir == 8'h1F)|(curr_ir == 8'h19)|(curr_ir == 8'hDF)|(curr_ir == 8'h1E)|(curr_ir == 8'hFE)|(curr_ir == 8'h07)|(curr_ir == 8'h5E)|(curr_ir == 8'h5F)|(curr_ir == 8'h1D)|(curr_ir == 8'h5D)|(curr_ir == 8'h1B)|(curr_ir == 8'hDD)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h46)|(curr_ir == 8'h06)|(curr_ir == 8'hC4)|(curr_ir == 8'h47)|(curr_ir == 8'h45)|(curr_ir == 8'h25)|(curr_ir == 8'hC5)|(curr_ir == 8'hE4)|(curr_ir == 8'h05)|(curr_ir == 8'hC7)|(curr_ir == 8'hE6)|(curr_ir == 8'hC6)|(curr_ir == 8'h07)|(curr_ir == 8'h24)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h33)|(curr_ir == 8'h43)|(curr_ir == 8'h13)|(curr_ir == 8'h03)|(curr_ir == 8'h53)|(curr_ir == 8'h23)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hC0)|(curr_ir == 8'h49)|(curr_ir == 8'hC9)|(curr_ir == 8'h4A)|(curr_ir == 8'h09)|(curr_ir == 8'hE0)|(curr_ir == 8'h0A)|(curr_ir == 8'h29)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h1F)|(curr_ir == 8'h3F)|(curr_ir == 8'h5B)|(curr_ir == 8'h1B)|(curr_ir == 8'h3B)|(curr_ir == 8'h5F))))
		alu_in_c = 0;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h0F)|(curr_ir == 8'h57)|(curr_ir == 8'h01)|(curr_ir == 8'h83)|(curr_ir == 8'hF1)|(curr_ir == 8'hD3)|(curr_ir == 8'h31)|(curr_ir == 8'h2F)|(curr_ir == 8'h41)|(curr_ir == 8'hE1)|(curr_ir == 8'hC1)|(curr_ir == 8'h71)|(curr_ir == 8'h37)|(curr_ir == 8'hF3)|(curr_ir == 8'hE3)|(curr_ir == 8'hD1)|(curr_ir == 8'h6F)|(curr_ir == 8'hC3)|(curr_ir == 8'h21)|(curr_ir == 8'h17)|(curr_ir == 8'h11)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h4F)|(curr_ir == 8'h77)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hF7)|(curr_ir == 8'hED)|(curr_ir == 8'hF5)|(curr_ir == 8'h35)|(curr_ir == 8'hEF)|(curr_ir == 8'h97)|(curr_ir == 8'h75)|(curr_ir == 8'h2D)|(curr_ir == 8'hCD)|(curr_ir == 8'hD5)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'h8F)|(curr_ir == 8'hD7)|(curr_ir == 8'h4D)|(curr_ir == 8'h6D)|(curr_ir == 8'hCF)|(curr_ir == 8'h0D)|(curr_ir == 8'h2C)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hD9)|(curr_ir == 8'hDB)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'h27)|(curr_ir == 8'hF9)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'hFF)|(curr_ir == 8'h19)|(curr_ir == 8'hDF)|(curr_ir == 8'h79)|(curr_ir == 8'h07)|(curr_ir == 8'h7D)|(curr_ir == 8'h1D)|(curr_ir == 8'hFB)|(curr_ir == 8'h67)|(curr_ir == 8'h5D)|(curr_ir == 8'hDD)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h33)|(curr_ir == 8'h73)|(curr_ir == 8'h63)|(curr_ir == 8'h43)|(curr_ir == 8'h13)|(curr_ir == 8'h03)|(curr_ir == 8'h53)|(curr_ir == 8'h23)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h1F)|(curr_ir == 8'h3F)|(curr_ir == 8'h5B)|(curr_ir == 8'h1B)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h7F)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h49)|(curr_ir == 8'hC9)|(curr_ir == 8'h4A)|(curr_ir == 8'h09)|(curr_ir == 8'hEB)|(curr_ir == 8'h69)|(curr_ir == 8'h6A)|(curr_ir == 8'hCB)|(curr_ir == 8'h2A)|(curr_ir == 8'hE9)|(curr_ir == 8'h0A)|(curr_ir == 8'h29)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h87)|(curr_ir == 8'hE7)|(curr_ir == 8'h45)|(curr_ir == 8'h25)|(curr_ir == 8'h65)|(curr_ir == 8'hC5)|(curr_ir == 8'hE5)|(curr_ir == 8'h05)|(curr_ir == 8'hC7)|(curr_ir == 8'h24))))
		alu_in_lhs = curr_a;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h0F)|(curr_ir == 8'h57)|(curr_ir == 8'h01)|(curr_ir == 8'hF1)|(curr_ir == 8'h31)|(curr_ir == 8'h2F)|(curr_ir == 8'h41)|(curr_ir == 8'hE1)|(curr_ir == 8'hC1)|(curr_ir == 8'h71)|(curr_ir == 8'h37)|(curr_ir == 8'hD1)|(curr_ir == 8'h6F)|(curr_ir == 8'h21)|(curr_ir == 8'h17)|(curr_ir == 8'h11)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h4F)|(curr_ir == 8'h77)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hED)|(curr_ir == 8'hF5)|(curr_ir == 8'h35)|(curr_ir == 8'h75)|(curr_ir == 8'h2D)|(curr_ir == 8'hCC)|(curr_ir == 8'hCD)|(curr_ir == 8'hD5)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'h4D)|(curr_ir == 8'h6D)|(curr_ir == 8'hEC)|(curr_ir == 8'h0D)|(curr_ir == 8'h2C)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hD9)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'h27)|(curr_ir == 8'hF9)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'h19)|(curr_ir == 8'h79)|(curr_ir == 8'h07)|(curr_ir == 8'h7D)|(curr_ir == 8'h1D)|(curr_ir == 8'h67)|(curr_ir == 8'h5D)|(curr_ir == 8'hDD)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h33)|(curr_ir == 8'h73)|(curr_ir == 8'h63)|(curr_ir == 8'h43)|(curr_ir == 8'h13)|(curr_ir == 8'h03)|(curr_ir == 8'h53)|(curr_ir == 8'h23)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hC0)|(curr_ir == 8'h49)|(curr_ir == 8'hC9)|(curr_ir == 8'h09)|(curr_ir == 8'hEB)|(curr_ir == 8'h69)|(curr_ir == 8'hE0)|(curr_ir == 8'hE9)|(curr_ir == 8'h29)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h1F)|(curr_ir == 8'h3F)|(curr_ir == 8'h5B)|(curr_ir == 8'h1B)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h7F)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hC4)|(curr_ir == 8'h45)|(curr_ir == 8'h25)|(curr_ir == 8'h65)|(curr_ir == 8'hC5)|(curr_ir == 8'hE5)|(curr_ir == 8'hE4)|(curr_ir == 8'h05)|(curr_ir == 8'h24))))
		alu_in_rhs = G_rd_data;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h0F)|(curr_ir == 8'h01)|(curr_ir == 8'h17)|(curr_ir == 8'h11)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h1F)|(curr_ir == 8'h1B)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h13)|(curr_ir == 8'h03)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h19)|(curr_ir == 8'h07)|(curr_ir == 8'h1D)))|
	    ((curr_cycle == 1)&(curr_ir == 8'h09))|
	    ((curr_cycle == 3)&((curr_ir == 8'h0D)|(curr_ir == 8'h15)))|
	    ((curr_cycle == 2)&(curr_ir == 8'h05)))
		next_a = alu_or;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h0F)|(curr_ir == 8'h57)|(curr_ir == 8'h01)|(curr_ir == 8'hA1)|(curr_ir == 8'hF1)|(curr_ir == 8'hEF)|(curr_ir == 8'h31)|(curr_ir == 8'h41)|(curr_ir == 8'hE1)|(curr_ir == 8'h71)|(curr_ir == 8'hF7)|(curr_ir == 8'h6F)|(curr_ir == 8'hB1)|(curr_ir == 8'h21)|(curr_ir == 8'h17)|(curr_ir == 8'h11)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h4F)|(curr_ir == 8'h77)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hED)|(curr_ir == 8'hF5)|(curr_ir == 8'h35)|(curr_ir == 8'h75)|(curr_ir == 8'h2D)|(curr_ir == 8'hAD)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'hB5)|(curr_ir == 8'h4D)|(curr_ir == 8'h6D)|(curr_ir == 8'h0D)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hE7)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'hF9)|(curr_ir == 8'hB9)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'h19)|(curr_ir == 8'h79)|(curr_ir == 8'h07)|(curr_ir == 8'h7D)|(curr_ir == 8'hBD)|(curr_ir == 8'h1D)|(curr_ir == 8'h67)|(curr_ir == 8'h5D)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hFF)|(curr_ir == 8'h1F)|(curr_ir == 8'hFB)|(curr_ir == 8'h5B)|(curr_ir == 8'h1B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h7F)))|
	    ((curr_cycle == 7)&((curr_ir == 8'hE3)|(curr_ir == 8'h73)|(curr_ir == 8'h63)|(curr_ir == 8'h43)|(curr_ir == 8'h13)|(curr_ir == 8'hF3)|(curr_ir == 8'h03)|(curr_ir == 8'h53)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h49)|(curr_ir == 8'h4A)|(curr_ir == 8'h09)|(curr_ir == 8'hEB)|(curr_ir == 8'h69)|(curr_ir == 8'hA9)|(curr_ir == 8'h6A)|(curr_ir == 8'h98)|(curr_ir == 8'h2A)|(curr_ir == 8'hE9)|(curr_ir == 8'h0A)|(curr_ir == 8'h29)|(curr_ir == 8'h8A)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hA5)|(curr_ir == 8'h45)|(curr_ir == 8'h25)|(curr_ir == 8'h65)|(curr_ir == 8'hE5)|(curr_ir == 8'h05))))
		next_p[Z_bit] = next_a == 0;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h0F)|(curr_ir == 8'h57)|(curr_ir == 8'h01)|(curr_ir == 8'hA1)|(curr_ir == 8'hF1)|(curr_ir == 8'hEF)|(curr_ir == 8'h31)|(curr_ir == 8'h41)|(curr_ir == 8'hE1)|(curr_ir == 8'h71)|(curr_ir == 8'hF7)|(curr_ir == 8'h6F)|(curr_ir == 8'hB1)|(curr_ir == 8'h21)|(curr_ir == 8'h17)|(curr_ir == 8'h11)|(curr_ir == 8'h61)|(curr_ir == 8'h51)|(curr_ir == 8'h4F)|(curr_ir == 8'h77)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hED)|(curr_ir == 8'hF5)|(curr_ir == 8'h35)|(curr_ir == 8'h75)|(curr_ir == 8'h2D)|(curr_ir == 8'hAD)|(curr_ir == 8'h15)|(curr_ir == 8'h55)|(curr_ir == 8'hB5)|(curr_ir == 8'h4D)|(curr_ir == 8'h6D)|(curr_ir == 8'h0D)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hE7)|(curr_ir == 8'h39)|(curr_ir == 8'hFD)|(curr_ir == 8'hF9)|(curr_ir == 8'hB9)|(curr_ir == 8'h59)|(curr_ir == 8'h3D)|(curr_ir == 8'h19)|(curr_ir == 8'h79)|(curr_ir == 8'h07)|(curr_ir == 8'h7D)|(curr_ir == 8'hBD)|(curr_ir == 8'h1D)|(curr_ir == 8'h67)|(curr_ir == 8'h5D)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hFF)|(curr_ir == 8'h1F)|(curr_ir == 8'hFB)|(curr_ir == 8'h5B)|(curr_ir == 8'h1B)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h7F)))|
	    ((curr_cycle == 7)&((curr_ir == 8'hE3)|(curr_ir == 8'h73)|(curr_ir == 8'h63)|(curr_ir == 8'h43)|(curr_ir == 8'h13)|(curr_ir == 8'hF3)|(curr_ir == 8'h03)|(curr_ir == 8'h53)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h49)|(curr_ir == 8'h4A)|(curr_ir == 8'h09)|(curr_ir == 8'hEB)|(curr_ir == 8'h69)|(curr_ir == 8'hA9)|(curr_ir == 8'h6A)|(curr_ir == 8'h98)|(curr_ir == 8'h2A)|(curr_ir == 8'hE9)|(curr_ir == 8'h0A)|(curr_ir == 8'h29)|(curr_ir == 8'h8A)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hA5)|(curr_ir == 8'h45)|(curr_ir == 8'h25)|(curr_ir == 8'h65)|(curr_ir == 8'hE5)|(curr_ir == 8'h05))))
		next_p[N_bit] = next_a[7];
	
	if (((curr_cycle == 1)&((curr_ir == 8'h22)|(curr_ir == 8'h52)|(curr_ir == 8'h82)|(curr_ir == 8'h42)|(curr_ir == 8'h02)|(curr_ir == 8'hB2)|(curr_ir == 8'hD2)|(curr_ir == 8'h32)|(curr_ir == 8'h92)|(curr_ir == 8'hF2)|(curr_ir == 8'h72)|(curr_ir == 8'h62)|(curr_ir == 8'h12))))
		next_cycle = -1;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h0F)|(curr_ir == 8'h76)|(curr_ir == 8'h37)|(curr_ir == 8'hD6)|(curr_ir == 8'h2E)|(curr_ir == 8'h0E)|(curr_ir == 8'h57)|(curr_ir == 8'h56)|(curr_ir == 8'hF6)|(curr_ir == 8'h6E)|(curr_ir == 8'h6F)|(curr_ir == 8'h16)|(curr_ir == 8'h4F)|(curr_ir == 8'h17)|(curr_ir == 8'h77)|(curr_ir == 8'h2F)|(curr_ir == 8'hEE)|(curr_ir == 8'hCE)|(curr_ir == 8'h36)|(curr_ir == 8'h4E)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h03)|(curr_ir == 8'h73)|(curr_ir == 8'h33)|(curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'h43)|(curr_ir == 8'h23)|(curr_ir == 8'h13)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h5F)|(curr_ir == 8'hDE)|(curr_ir == 8'hFE)|(curr_ir == 8'h5B)|(curr_ir == 8'h5E)|(curr_ir == 8'h1F)|(curr_ir == 8'h1B)|(curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h1E)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h46)|(curr_ir == 8'h67)|(curr_ir == 8'h06)|(curr_ir == 8'h07)|(curr_ir == 8'h26)|(curr_ir == 8'h27)|(curr_ir == 8'h66)|(curr_ir == 8'hE6)|(curr_ir == 8'h47)|(curr_ir == 8'hC6))))
		alu_in_lhs = G_rd_data;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h0F)|(curr_ir == 8'h76)|(curr_ir == 8'h37)|(curr_ir == 8'h2E)|(curr_ir == 8'h0E)|(curr_ir == 8'h57)|(curr_ir == 8'h56)|(curr_ir == 8'h6E)|(curr_ir == 8'h6F)|(curr_ir == 8'h16)|(curr_ir == 8'h4F)|(curr_ir == 8'h17)|(curr_ir == 8'h77)|(curr_ir == 8'h2F)|(curr_ir == 8'h36)|(curr_ir == 8'h4E)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h03)|(curr_ir == 8'h73)|(curr_ir == 8'h33)|(curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'h43)|(curr_ir == 8'h23)|(curr_ir == 8'h13)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h5F)|(curr_ir == 8'h5B)|(curr_ir == 8'h5E)|(curr_ir == 8'h1F)|(curr_ir == 8'h1B)|(curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h1E)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h4A)|(curr_ir == 8'h0A)|(curr_ir == 8'h2A)|(curr_ir == 8'h6A)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h46)|(curr_ir == 8'h67)|(curr_ir == 8'h06)|(curr_ir == 8'h07)|(curr_ir == 8'h26)|(curr_ir == 8'h27)|(curr_ir == 8'h66)|(curr_ir == 8'h47))))
		alu_in_rhs = 0;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h26)|(curr_ir == 8'h27)|(curr_ir == 8'h07)|(curr_ir == 8'h06)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h1B)|(curr_ir == 8'h1E)|(curr_ir == 8'h3E)|(curr_ir == 8'h3F)|(curr_ir == 8'h2E)|(curr_ir == 8'h0E)|(curr_ir == 8'h3B)|(curr_ir == 8'h16)|(curr_ir == 8'h36)|(curr_ir == 8'h1F)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h17)|(curr_ir == 8'h16)|(curr_ir == 8'h2F)|(curr_ir == 8'h06)|(curr_ir == 8'h36)|(curr_ir == 8'h26)|(curr_ir == 8'h37)|(curr_ir == 8'h0F)|(curr_ir == 8'h2E)|(curr_ir == 8'h0E)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'h03)|(curr_ir == 8'h33)|(curr_ir == 8'h1E)|(curr_ir == 8'h3E))))
		G_wr_data = alu_rol;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h27)|(curr_ir == 8'h07)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h1B)|(curr_ir == 8'h3F)|(curr_ir == 8'h2E)|(curr_ir == 8'h0E)|(curr_ir == 8'h3B)|(curr_ir == 8'h16)|(curr_ir == 8'h36)|(curr_ir == 8'h1F)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h17)|(curr_ir == 8'h2F)|(curr_ir == 8'h06)|(curr_ir == 8'h26)|(curr_ir == 8'h37)|(curr_ir == 8'h0F)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h23)|(curr_ir == 8'h13)|(curr_ir == 8'h03)|(curr_ir == 8'h33)|(curr_ir == 8'h1E)|(curr_ir == 8'h3E)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h0A)|(curr_ir == 8'h2A))))
		next_p[C_bit] = alu_rol_c;
	
	if (((curr_cycle == 1)&((curr_ir == 8'hD1)|(curr_ir == 8'hD7)|(curr_ir == 8'hC7)|(curr_ir == 8'hF5)|(curr_ir == 8'h34)|(curr_ir == 8'h95)|(curr_ir == 8'h85)|(curr_ir == 8'hC5)|(curr_ir == 8'h86)|(curr_ir == 8'h14)|(curr_ir == 8'h65)|(curr_ir == 8'hC6)|(curr_ir == 8'h17)|(curr_ir == 8'h11)|(curr_ir == 8'h53)|(curr_ir == 8'hB4)|(curr_ir == 8'h77)|(curr_ir == 8'h67)|(curr_ir == 8'h84)|(curr_ir == 8'h35)|(curr_ir == 8'h66)|(curr_ir == 8'h54)|(curr_ir == 8'h73)|(curr_ir == 8'h33)|(curr_ir == 8'h57)|(curr_ir == 8'h94)|(curr_ir == 8'h25)|(curr_ir == 8'hE6)|(curr_ir == 8'h55)|(curr_ir == 8'hB6)|(curr_ir == 8'h07)|(curr_ir == 8'h06)|(curr_ir == 8'hE4)|(curr_ir == 8'hF1)|(curr_ir == 8'hD5)|(curr_ir == 8'h26)|(curr_ir == 8'h37)|(curr_ir == 8'h05)|(curr_ir == 8'hA5)|(curr_ir == 8'hD3)|(curr_ir == 8'h24)|(curr_ir == 8'h31)|(curr_ir == 8'hB7)|(curr_ir == 8'hC4)|(curr_ir == 8'h15)|(curr_ir == 8'h91)|(curr_ir == 8'h97)|(curr_ir == 8'h87)|(curr_ir == 8'h75)|(curr_ir == 8'hB5)|(curr_ir == 8'h13)|(curr_ir == 8'hA6)|(curr_ir == 8'hD4)|(curr_ir == 8'h76)|(curr_ir == 8'h74)|(curr_ir == 8'h64)|(curr_ir == 8'h71)|(curr_ir == 8'hA4)|(curr_ir == 8'hB1)|(curr_ir == 8'h27)|(curr_ir == 8'h44)|(curr_ir == 8'hF6)|(curr_ir == 8'h47)|(curr_ir == 8'h56)|(curr_ir == 8'hA7)|(curr_ir == 8'hE7)|(curr_ir == 8'h16)|(curr_ir == 8'hF4)|(curr_ir == 8'h46)|(curr_ir == 8'hE5)|(curr_ir == 8'h36)|(curr_ir == 8'h51)|(curr_ir == 8'h45)|(curr_ir == 8'h96)|(curr_ir == 8'hF7)|(curr_ir == 8'hB3)|(curr_ir == 8'h04)|(curr_ir == 8'hD6)|(curr_ir == 8'hF3))))
		next_adh = 0;
	
	if (((curr_cycle == 4)&((curr_ir == 8'h2F)|(curr_ir == 8'h06)|(curr_ir == 8'h26)|(curr_ir == 8'h37)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h23)|(curr_ir == 8'h33)|(curr_ir == 8'h1E)|(curr_ir == 8'h3E)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h3F)|(curr_ir == 8'h16)|(curr_ir == 8'h36)|(curr_ir == 8'h2E)|(curr_ir == 8'h0E)|(curr_ir == 8'h3B)))|
	    ((curr_cycle == 3)&(curr_ir == 8'h27)))
		next_p[Z_bit] = alu_rol == 0;
	
	if (((curr_cycle == 4)&((curr_ir == 8'h2F)|(curr_ir == 8'h06)|(curr_ir == 8'h26)|(curr_ir == 8'h37)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h23)|(curr_ir == 8'h33)|(curr_ir == 8'h1E)|(curr_ir == 8'h3E)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h3F)|(curr_ir == 8'h16)|(curr_ir == 8'h36)|(curr_ir == 8'h2E)|(curr_ir == 8'h0E)|(curr_ir == 8'h3B)))|
	    ((curr_cycle == 3)&(curr_ir == 8'h27)))
		next_p[N_bit] = alu_rol[7];
	
	if (((curr_cycle == 2)&(curr_ir == 8'h08)))
		G_wr_data = curr_p | B_mask;
	
	if (((curr_cycle == 1)&((curr_ir == 8'h2A)|(curr_ir == 8'h0A))))
		next_a = alu_rol;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h0F)|(curr_ir == 8'hAE)|(curr_ir == 8'h8C)|(curr_ir == 8'hED)|(curr_ir == 8'h4D)|(curr_ir == 8'hAF)|(curr_ir == 8'hEF)|(curr_ir == 8'h2E)|(curr_ir == 8'h0C)|(curr_ir == 8'h6D)|(curr_ir == 8'h0E)|(curr_ir == 8'hCF)|(curr_ir == 8'hEC)|(curr_ir == 8'h6E)|(curr_ir == 8'hAD)|(curr_ir == 8'h6F)|(curr_ir == 8'h4F)|(curr_ir == 8'h2D)|(curr_ir == 8'hCC)|(curr_ir == 8'h8D)|(curr_ir == 8'h8E)|(curr_ir == 8'h2F)|(curr_ir == 8'hCD)|(curr_ir == 8'hEE)|(curr_ir == 8'hCE)|(curr_ir == 8'hAC)|(curr_ir == 8'h8F)|(curr_ir == 8'h2C)|(curr_ir == 8'h0D)|(curr_ir == 8'h4E))))
		{next_pch, next_pcl} = curr_pc;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h10)))
		next_cycle = (curr_p[N_bit] ? 0 : (curr_cycle + 1));
	
	if (((curr_cycle == 1)&((curr_ir == 8'h70)|(curr_ir == 8'h30)|(curr_ir == 8'h50)|(curr_ir == 8'h10)|(curr_ir == 8'hB0)|(curr_ir == 8'hD0)|(curr_ir == 8'h90)|(curr_ir == 8'hF0))))
		{next_adh, next_adl} = {8'h00, G_rd_data} + (curr_pc + 1) - {7'h00, G_rd_data[7], 8'h00};
	
	if (((curr_cycle == 2)&((curr_ir == 8'h10)|(curr_ir == 8'hD0)|(curr_ir == 8'h30)|(curr_ir == 8'h50)|(curr_ir == 8'hF0)|(curr_ir == 8'hB0)|(curr_ir == 8'h70)|(curr_ir == 8'h90))))
		G_addr = {curr_pch, curr_adl};
	
	if (((curr_cycle == 2)&((curr_ir == 8'h10)|(curr_ir == 8'hD0)|(curr_ir == 8'h30)|(curr_ir == 8'h50)|(curr_ir == 8'hF0)|(curr_ir == 8'hB0)|(curr_ir == 8'h70)|(curr_ir == 8'h90))))
		{next_pch, next_pcl} = curr_ad;
	
	if (((curr_cycle == 2)&((curr_ir == 8'h10)|(curr_ir == 8'hD0)|(curr_ir == 8'h30)|(curr_ir == 8'h50)|(curr_ir == 8'hF0)|(curr_ir == 8'hB0)|(curr_ir == 8'h70)|(curr_ir == 8'h90))))
		next_cycle = ((curr_adh != curr_pch) ? (curr_cycle + 1) : 0);
	
	if (((curr_cycle == 2)&((curr_ir == 8'h71)|(curr_ir == 8'hB3)|(curr_ir == 8'h13)|(curr_ir == 8'hD1)|(curr_ir == 8'h91)|(curr_ir == 8'hB1)|(curr_ir == 8'h33)|(curr_ir == 8'hD3)|(curr_ir == 8'hF3)|(curr_ir == 8'h11)|(curr_ir == 8'h53)|(curr_ir == 8'h31)|(curr_ir == 8'h73)|(curr_ir == 8'h51)|(curr_ir == 8'hF1))))
		next_adl = curr_adl + 1;
	
	if (((curr_cycle == 2)&((curr_ir == 8'hFF)|(curr_ir == 8'h5F)|(curr_ir == 8'h39)|(curr_ir == 8'h6C)|(curr_ir == 8'hFE)|(curr_ir == 8'h5C)|(curr_ir == 8'hFB)|(curr_ir == 8'hD9)|(curr_ir == 8'hBC)|(curr_ir == 8'h5B)|(curr_ir == 8'h5E)|(curr_ir == 8'hDE)|(curr_ir == 8'h1D)|(curr_ir == 8'h1F)|(curr_ir == 8'hBE)|(curr_ir == 8'h5D)|(curr_ir == 8'hFC)|(curr_ir == 8'hBF)|(curr_ir == 8'h99)|(curr_ir == 8'h1B)|(curr_ir == 8'hFD)|(curr_ir == 8'h1C)|(curr_ir == 8'h3F)|(curr_ir == 8'h7C)|(curr_ir == 8'h7D)|(curr_ir == 8'h1E)|(curr_ir == 8'h7F)|(curr_ir == 8'h3E)|(curr_ir == 8'hDD)|(curr_ir == 8'hF9)|(curr_ir == 8'hBD)|(curr_ir == 8'h3B)|(curr_ir == 8'h7E)|(curr_ir == 8'hDB)|(curr_ir == 8'h19)|(curr_ir == 8'h7B)|(curr_ir == 8'h59)|(curr_ir == 8'hDF)|(curr_ir == 8'h79)|(curr_ir == 8'hB9)|(curr_ir == 8'h3D)|(curr_ir == 8'h9D)|(curr_ir == 8'hDC)|(curr_ir == 8'h3C)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h71)|(curr_ir == 8'h73)|(curr_ir == 8'hD1)|(curr_ir == 8'hD3)|(curr_ir == 8'hB1)|(curr_ir == 8'h33)|(curr_ir == 8'h53)|(curr_ir == 8'h31)|(curr_ir == 8'h91)|(curr_ir == 8'h11)|(curr_ir == 8'h13)|(curr_ir == 8'hF1)|(curr_ir == 8'h51)|(curr_ir == 8'hF3)|(curr_ir == 8'hB3))))
		next_bah = G_rd_data;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h71)|(curr_ir == 8'h73)|(curr_ir == 8'hD1)|(curr_ir == 8'hD3)|(curr_ir == 8'hB1)|(curr_ir == 8'h33)|(curr_ir == 8'h53)|(curr_ir == 8'h31)|(curr_ir == 8'h91)|(curr_ir == 8'h11)|(curr_ir == 8'h13)|(curr_ir == 8'hF1)|(curr_ir == 8'h51)|(curr_ir == 8'hF3)|(curr_ir == 8'hB3)))|
	    ((curr_cycle == 2)&((curr_ir == 8'h39)|(curr_ir == 8'hFB)|(curr_ir == 8'hD9)|(curr_ir == 8'h5B)|(curr_ir == 8'hBE)|(curr_ir == 8'hBF)|(curr_ir == 8'h99)|(curr_ir == 8'h1B)|(curr_ir == 8'hF9)|(curr_ir == 8'h3B)|(curr_ir == 8'h19)|(curr_ir == 8'h7B)|(curr_ir == 8'h59)|(curr_ir == 8'h79)|(curr_ir == 8'hB9)|(curr_ir == 8'hDB))))
		{next_adh, next_adl} = {G_rd_data, curr_bal}  + {8'h00, curr_y};
	
	if (((curr_cycle == 2)&((curr_ir == 8'hFF)|(curr_ir == 8'h5F)|(curr_ir == 8'h39)|(curr_ir == 8'h5C)|(curr_ir == 8'hFB)|(curr_ir == 8'hD9)|(curr_ir == 8'hBC)|(curr_ir == 8'h5B)|(curr_ir == 8'h1D)|(curr_ir == 8'h1F)|(curr_ir == 8'hBE)|(curr_ir == 8'h5D)|(curr_ir == 8'hFC)|(curr_ir == 8'hBF)|(curr_ir == 8'h1B)|(curr_ir == 8'hFD)|(curr_ir == 8'h1C)|(curr_ir == 8'h3F)|(curr_ir == 8'h7C)|(curr_ir == 8'h7D)|(curr_ir == 8'h7F)|(curr_ir == 8'hF9)|(curr_ir == 8'hDD)|(curr_ir == 8'hBD)|(curr_ir == 8'h3B)|(curr_ir == 8'hDB)|(curr_ir == 8'h19)|(curr_ir == 8'h7B)|(curr_ir == 8'h59)|(curr_ir == 8'hDF)|(curr_ir == 8'h79)|(curr_ir == 8'hB9)|(curr_ir == 8'h3D)|(curr_ir == 8'hDC)|(curr_ir == 8'h3C)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h71)|(curr_ir == 8'h73)|(curr_ir == 8'hD1)|(curr_ir == 8'hD3)|(curr_ir == 8'hB1)|(curr_ir == 8'h33)|(curr_ir == 8'h53)|(curr_ir == 8'h31)|(curr_ir == 8'h11)|(curr_ir == 8'h13)|(curr_ir == 8'hF1)|(curr_ir == 8'h51)|(curr_ir == 8'hF3)|(curr_ir == 8'hB3))))
		next_cycle = curr_cycle + 1 + ((next_bah != next_adh) ? 0 : 1);
	
	if (((curr_cycle == 3)&((curr_ir == 8'h3E)|(curr_ir == 8'hBE)|(curr_ir == 8'h7D)|(curr_ir == 8'hBF)|(curr_ir == 8'h1C)|(curr_ir == 8'h99)|(curr_ir == 8'h3F)|(curr_ir == 8'h1E)|(curr_ir == 8'hF9)|(curr_ir == 8'hDD)|(curr_ir == 8'h7E)|(curr_ir == 8'hBD)|(curr_ir == 8'h7C)|(curr_ir == 8'h3B)|(curr_ir == 8'h19)|(curr_ir == 8'h7F)|(curr_ir == 8'h59)|(curr_ir == 8'h79)|(curr_ir == 8'hB9)|(curr_ir == 8'hDF)|(curr_ir == 8'h5F)|(curr_ir == 8'h3D)|(curr_ir == 8'h7B)|(curr_ir == 8'h3C)|(curr_ir == 8'hDB)|(curr_ir == 8'h39)|(curr_ir == 8'h9D)|(curr_ir == 8'hDE)|(curr_ir == 8'hFE)|(curr_ir == 8'hDC)|(curr_ir == 8'h1D)|(curr_ir == 8'hFF)|(curr_ir == 8'h5C)|(curr_ir == 8'hD9)|(curr_ir == 8'h5E)|(curr_ir == 8'h1F)|(curr_ir == 8'hFB)|(curr_ir == 8'hBC)|(curr_ir == 8'h5D)|(curr_ir == 8'h5B)|(curr_ir == 8'hFC)|(curr_ir == 8'h1B)|(curr_ir == 8'hFD)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h53)|(curr_ir == 8'h13)|(curr_ir == 8'h11)|(curr_ir == 8'h51)|(curr_ir == 8'hF1)|(curr_ir == 8'hB3)|(curr_ir == 8'hF3)|(curr_ir == 8'hD1)|(curr_ir == 8'h71)|(curr_ir == 8'hD3)|(curr_ir == 8'hB1)|(curr_ir == 8'h33)|(curr_ir == 8'h73)|(curr_ir == 8'h31)|(curr_ir == 8'h91))))
		G_addr = {curr_bah, curr_adl};
	
	if (((curr_cycle == 2)&((curr_ir == 8'h75)|(curr_ir == 8'h16)|(curr_ir == 8'hB4)|(curr_ir == 8'h55)|(curr_ir == 8'h17)|(curr_ir == 8'h77)|(curr_ir == 8'hB5)|(curr_ir == 8'h74)|(curr_ir == 8'hF4)|(curr_ir == 8'h35)|(curr_ir == 8'h36)|(curr_ir == 8'hD5)|(curr_ir == 8'h76)|(curr_ir == 8'h37)|(curr_ir == 8'hD4)|(curr_ir == 8'hF7)|(curr_ir == 8'hD7)|(curr_ir == 8'hD6)|(curr_ir == 8'h56)|(curr_ir == 8'h34)|(curr_ir == 8'h95)|(curr_ir == 8'h54)|(curr_ir == 8'h94)|(curr_ir == 8'h57)|(curr_ir == 8'hF6)|(curr_ir == 8'hF5)|(curr_ir == 8'h14)|(curr_ir == 8'h15))))
		next_adl = curr_adl + curr_x;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h18)))
		next_p[C_bit] = 0;
	
	if (((curr_cycle == 2)&((curr_ir == 8'hFF)|(curr_ir == 8'h5F)|(curr_ir == 8'hFE)|(curr_ir == 8'h5C)|(curr_ir == 8'hBC)|(curr_ir == 8'h5E)|(curr_ir == 8'hDE)|(curr_ir == 8'h1D)|(curr_ir == 8'h1F)|(curr_ir == 8'h5D)|(curr_ir == 8'hFC)|(curr_ir == 8'hFD)|(curr_ir == 8'h1C)|(curr_ir == 8'h3F)|(curr_ir == 8'h7C)|(curr_ir == 8'h7D)|(curr_ir == 8'h1E)|(curr_ir == 8'h7F)|(curr_ir == 8'h3E)|(curr_ir == 8'hDD)|(curr_ir == 8'hBD)|(curr_ir == 8'h7E)|(curr_ir == 8'hDF)|(curr_ir == 8'h3D)|(curr_ir == 8'h9D)|(curr_ir == 8'hDC)|(curr_ir == 8'h3C))))
		{next_adh, next_adl} = {G_rd_data, curr_bal}  + {8'h00, curr_x};
	
	if (((curr_cycle == 2)&(curr_ir == 8'h25))|
	    ((curr_cycle == 5)&((curr_ir == 8'h2F)|(curr_ir == 8'h37)|(curr_ir == 8'h21)|(curr_ir == 8'h31)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h35)|(curr_ir == 8'h2D)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h39)|(curr_ir == 8'h3D)|(curr_ir == 8'h27)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h23)|(curr_ir == 8'h33)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h3B)|(curr_ir == 8'h3F)))|
	    ((curr_cycle == 1)&(curr_ir == 8'h29)))
		next_a = alu_and;
	
	if (((curr_cycle == 5)&((curr_ir == 8'hF1)|(curr_ir == 8'h71)|(curr_ir == 8'hE1)|(curr_ir == 8'hF3)|(curr_ir == 8'hE3)|(curr_ir == 8'h73)|(curr_ir == 8'h33)|(curr_ir == 8'h63)|(curr_ir == 8'h6F)|(curr_ir == 8'h61)|(curr_ir == 8'h23)|(curr_ir == 8'h77)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hF7)|(curr_ir == 8'hED)|(curr_ir == 8'h76)|(curr_ir == 8'h37)|(curr_ir == 8'hEF)|(curr_ir == 8'h2E)|(curr_ir == 8'h6D)|(curr_ir == 8'hF5)|(curr_ir == 8'h6E)|(curr_ir == 8'h6F)|(curr_ir == 8'h75)|(curr_ir == 8'h77)|(curr_ir == 8'h2F)|(curr_ir == 8'h36)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hE7)|(curr_ir == 8'h67)|(curr_ir == 8'hE5)|(curr_ir == 8'h26)|(curr_ir == 8'h27)|(curr_ir == 8'h66)|(curr_ir == 8'h65)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hE9)|(curr_ir == 8'hEB)|(curr_ir == 8'h69)|(curr_ir == 8'h2A)|(curr_ir == 8'h6A)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h7B)|(curr_ir == 8'h7F)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hFF)|(curr_ir == 8'hFB)|(curr_ir == 8'hFD)|(curr_ir == 8'h67)|(curr_ir == 8'h7D)|(curr_ir == 8'hF9)|(curr_ir == 8'h3E)|(curr_ir == 8'h7E)|(curr_ir == 8'h3F)|(curr_ir == 8'h7F)|(curr_ir == 8'h79)|(curr_ir == 8'h3B)|(curr_ir == 8'h7B)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h73)|(curr_ir == 8'h63))))
		alu_in_c = curr_p[C_bit];
	
	if (((curr_cycle == 2)&(curr_ir == 8'h24))|
	    ((curr_cycle == 3)&(curr_ir == 8'h2C)))
		next_p[Z_bit] = alu_and == 0;
	
	if (((curr_cycle == 2)&(curr_ir == 8'h24))|
	    ((curr_cycle == 3)&(curr_ir == 8'h2C)))
		next_p[V_bit] = G_rd_data[6];
	
	if (((curr_cycle == 3)&((curr_ir == 8'h68)|(curr_ir == 8'h2C)))|
	    ((curr_cycle == 2)&(curr_ir == 8'h24)))
		next_p[N_bit] = G_rd_data[7];
	
	if (((curr_cycle == 2)&((curr_ir == 8'h68)|(curr_ir == 8'h40)|(curr_ir == 8'h60)|(curr_ir == 8'h28)))|
	    ((curr_cycle == 4)&(curr_ir == 8'h40))|
	    ((curr_cycle == 3)&((curr_ir == 8'h60)|(curr_ir == 8'h40))))
		next_s = curr_s + 1;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h28)|(curr_ir == 8'h40))))
		next_p = G_rd_data;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h30)))
		next_cycle = (curr_p[N_bit] ? (curr_cycle + 1) : 0);
	
	if (((curr_cycle == 1)&(curr_ir == 8'h38)))
		next_p[C_bit] = 1;
	
	if (((curr_cycle == 4)&(curr_ir == 8'h40))|
	    ((curr_cycle == 3)&(curr_ir == 8'h60)))
		next_pcl = G_rd_data;
	
	if (((curr_cycle == 5)&(curr_ir == 8'h40))|
	    ((curr_cycle == 4)&(curr_ir == 8'h60)))
		next_pch = G_rd_data;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h51)|(curr_ir == 8'h4F)|(curr_ir == 8'h41)|(curr_ir == 8'h57)))|
	    ((curr_cycle == 1)&(curr_ir == 8'h49))|
	    ((curr_cycle == 4)&((curr_ir == 8'h59)|(curr_ir == 8'h5D)|(curr_ir == 8'h47)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h4D)|(curr_ir == 8'h55)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h43)|(curr_ir == 8'h53)))|
	    ((curr_cycle == 2)&(curr_ir == 8'h45))|
	    ((curr_cycle == 6)&((curr_ir == 8'h5B)|(curr_ir == 8'h5F))))
		next_a = alu_xor;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h4E)|(curr_ir == 8'h56)|(curr_ir == 8'h7F)|(curr_ir == 8'h7E)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h6E)|(curr_ir == 8'h5B)|(curr_ir == 8'h5E)|(curr_ir == 8'h76)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h6F)|(curr_ir == 8'h77)|(curr_ir == 8'h4F)|(curr_ir == 8'h46)|(curr_ir == 8'h76)|(curr_ir == 8'h4E)|(curr_ir == 8'h66)|(curr_ir == 8'h56)|(curr_ir == 8'h57)|(curr_ir == 8'h6E)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'h43)|(curr_ir == 8'h5E)|(curr_ir == 8'h73)|(curr_ir == 8'h7E)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h66)|(curr_ir == 8'h47)|(curr_ir == 8'h46)|(curr_ir == 8'h67))))
		G_wr_data = alu_ror;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h4E)|(curr_ir == 8'h56)|(curr_ir == 8'h7F)|(curr_ir == 8'h7B)|(curr_ir == 8'h5F)|(curr_ir == 8'h6E)|(curr_ir == 8'h5B)|(curr_ir == 8'h76)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h6F)|(curr_ir == 8'h77)|(curr_ir == 8'h4F)|(curr_ir == 8'h46)|(curr_ir == 8'h66)|(curr_ir == 8'h57)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h63)|(curr_ir == 8'h53)|(curr_ir == 8'h43)|(curr_ir == 8'h5E)|(curr_ir == 8'h73)|(curr_ir == 8'h7E)))|
	    ((curr_cycle == 1)&((curr_ir == 8'h4A)|(curr_ir == 8'h6A)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h47)|(curr_ir == 8'h67))))
		next_p[C_bit] = alu_ror_c;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h4E)|(curr_ir == 8'h56)|(curr_ir == 8'h6E)|(curr_ir == 8'h76)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h46)|(curr_ir == 8'h66)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h7E)|(curr_ir == 8'h5E))))
		next_p[Z_bit] = alu_ror == 0;
	
	if (((curr_cycle == 5)&((curr_ir == 8'h4E)|(curr_ir == 8'h56)|(curr_ir == 8'h6E)|(curr_ir == 8'h76)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h46)|(curr_ir == 8'h66)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h7E)|(curr_ir == 8'h5E))))
		next_p[N_bit] = alu_ror[7];
	
	if (((curr_cycle == 2)&((curr_ir == 8'h85)|(curr_ir == 8'h48)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h95)|(curr_ir == 8'h8D)))|
	    ((curr_cycle == 4)&((curr_ir == 8'h99)|(curr_ir == 8'h9D)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h91)|(curr_ir == 8'h81))))
		G_wr_data = curr_a;
	
	if (((curr_cycle == 1)&((curr_ir == 8'h4A)|(curr_ir == 8'h6A))))
		next_a = alu_ror;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h50)))
		next_cycle = (curr_p[V_bit] ? 0 : (curr_cycle + 1));
	
	if (((curr_cycle == 1)&(curr_ir == 8'h58)))
		next_p[I_bit] = 0;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h6D)|(curr_ir == 8'h75)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h71)|(curr_ir == 8'h77)|(curr_ir == 8'h6F)|(curr_ir == 8'h61)))|
	    ((curr_cycle == 2)&(curr_ir == 8'h65))|
	    ((curr_cycle == 4)&((curr_ir == 8'h67)|(curr_ir == 8'h79)|(curr_ir == 8'h7D)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h7F)|(curr_ir == 8'h7B)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h73)|(curr_ir == 8'h63)))|
	    ((curr_cycle == 1)&(curr_ir == 8'h69)))
		next_a = alu_adc[7:0];
	
	if (((curr_cycle == 3)&((curr_ir == 8'h6D)|(curr_ir == 8'h75)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h71)|(curr_ir == 8'h77)|(curr_ir == 8'h6F)|(curr_ir == 8'h61)))|
	    ((curr_cycle == 2)&(curr_ir == 8'h65))|
	    ((curr_cycle == 4)&((curr_ir == 8'h67)|(curr_ir == 8'h79)|(curr_ir == 8'h7D)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h7F)|(curr_ir == 8'h7B)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h73)|(curr_ir == 8'h63)))|
	    ((curr_cycle == 1)&(curr_ir == 8'h69)))
		next_p[C_bit] = alu_adc_c;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h6D)|(curr_ir == 8'h75)))|
	    ((curr_cycle == 5)&((curr_ir == 8'h71)|(curr_ir == 8'h77)|(curr_ir == 8'h6F)|(curr_ir == 8'h61)))|
	    ((curr_cycle == 2)&(curr_ir == 8'h65))|
	    ((curr_cycle == 4)&((curr_ir == 8'h67)|(curr_ir == 8'h79)|(curr_ir == 8'h7D)))|
	    ((curr_cycle == 6)&((curr_ir == 8'h7F)|(curr_ir == 8'h7B)))|
	    ((curr_cycle == 7)&((curr_ir == 8'h73)|(curr_ir == 8'h63)))|
	    ((curr_cycle == 1)&(curr_ir == 8'h69)))
		next_p[V_bit] = alu_adc_v;
	
	if (((curr_cycle == 4)&((curr_ir == 8'hBD)|(curr_ir == 8'hBF)|(curr_ir == 8'hB9)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hA9)|(curr_ir == 8'hAB)))|
	    ((curr_cycle == 3)&((curr_ir == 8'h68)|(curr_ir == 8'hAF)|(curr_ir == 8'hB7)|(curr_ir == 8'hAD)|(curr_ir == 8'hB5)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hA5)|(curr_ir == 8'hA7)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hA1)|(curr_ir == 8'hB1)|(curr_ir == 8'hB3)|(curr_ir == 8'hA3))))
		next_a = G_rd_data;
	
	if (((curr_cycle == 3)&(curr_ir == 8'h68)))
		next_p[Z_bit] = G_rd_data == 0;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h70)))
		next_cycle = (curr_p[V_bit] ? (curr_cycle + 1) : 0);
	
	if (((curr_cycle == 1)&(curr_ir == 8'h78)))
		next_p[I_bit] = 1;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h8F)|(curr_ir == 8'h97)))|
	    ((curr_cycle == 5)&(curr_ir == 8'h83))|
	    ((curr_cycle == 1)&(curr_ir == 8'hCB))|
	    ((curr_cycle == 2)&(curr_ir == 8'h87)))
		alu_in_rhs = curr_x;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h8F)|(curr_ir == 8'h97)))|
	    ((curr_cycle == 5)&(curr_ir == 8'h83))|
	    ((curr_cycle == 1)&(curr_ir == 8'hCB))|
	    ((curr_cycle == 2)&(curr_ir == 8'h87)))
		G_wr_data = alu_and;
	
	if (((curr_cycle == 2)&(curr_ir == 8'h84))|
	    ((curr_cycle == 3)&((curr_ir == 8'h8C)|(curr_ir == 8'h94))))
		G_wr_data = curr_y;
	
	if (((curr_cycle == 3)&((curr_ir == 8'h96)|(curr_ir == 8'h8E)))|
	    ((curr_cycle == 2)&(curr_ir == 8'h86)))
		G_wr_data = curr_x;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h88)))
		next_y = curr_y - 1;
	
	if (((curr_cycle == 2)&(curr_ir == 8'hA4))|
	    ((curr_cycle == 1)&((curr_ir == 8'hA8)|(curr_ir == 8'hC8)|(curr_ir == 8'hA0)|(curr_ir == 8'h88)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hAC)|(curr_ir == 8'hB4)))|
	    ((curr_cycle == 4)&(curr_ir == 8'hBC)))
		next_p[Z_bit] = next_y == 0;
	
	if (((curr_cycle == 2)&(curr_ir == 8'hA4))|
	    ((curr_cycle == 1)&((curr_ir == 8'hA8)|(curr_ir == 8'hC8)|(curr_ir == 8'hA0)|(curr_ir == 8'h88)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hAC)|(curr_ir == 8'hB4)))|
	    ((curr_cycle == 4)&(curr_ir == 8'hBC)))
		next_p[N_bit] = next_y[7];
	
	if (((curr_cycle == 1)&(curr_ir == 8'h8A)))
		next_a = curr_x;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h90)))
		next_cycle = (curr_p[C_bit] ? 0 : (curr_cycle + 1));
	
	if (((curr_cycle == 2)&((curr_ir == 8'hB6)|(curr_ir == 8'hB7)|(curr_ir == 8'h96)|(curr_ir == 8'h97))))
		next_adl = curr_adl + curr_y;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h98)))
		next_a = curr_y;
	
	if (((curr_cycle == 1)&(curr_ir == 8'h9A)))
		next_s = curr_x;
	
	if (((curr_cycle == 2)&(curr_ir == 8'hA4))|
	    ((curr_cycle == 3)&((curr_ir == 8'hAC)|(curr_ir == 8'hB4)))|
	    ((curr_cycle == 4)&(curr_ir == 8'hBC))|
	    ((curr_cycle == 1)&(curr_ir == 8'hA0)))
		next_y = G_rd_data;
	
	if (((curr_cycle == 3)&((curr_ir == 8'hAE)|(curr_ir == 8'hAF)|(curr_ir == 8'hB6)|(curr_ir == 8'hB7)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hBE)|(curr_ir == 8'hBF)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hA2)|(curr_ir == 8'hAB)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hA7)|(curr_ir == 8'hA6)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hB3)|(curr_ir == 8'hA3))))
		next_x = G_rd_data;
	
	if (((curr_cycle == 1)&((curr_ir == 8'hBA)|(curr_ir == 8'hE8)|(curr_ir == 8'hA2)|(curr_ir == 8'hCA)|(curr_ir == 8'hAA)|(curr_ir == 8'hAB)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hAE)|(curr_ir == 8'hAF)|(curr_ir == 8'hB6)|(curr_ir == 8'hB7)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hBE)|(curr_ir == 8'hBF)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hA7)|(curr_ir == 8'hA6)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hB3)|(curr_ir == 8'hA3))))
		next_p[N_bit] = next_x[7];
	
	if (((curr_cycle == 1)&((curr_ir == 8'hBA)|(curr_ir == 8'hE8)|(curr_ir == 8'hA2)|(curr_ir == 8'hCA)|(curr_ir == 8'hAA)|(curr_ir == 8'hAB)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hAE)|(curr_ir == 8'hAF)|(curr_ir == 8'hB6)|(curr_ir == 8'hB7)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hBE)|(curr_ir == 8'hBF)))|
	    ((curr_cycle == 2)&((curr_ir == 8'hA7)|(curr_ir == 8'hA6)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hB3)|(curr_ir == 8'hA3))))
		next_p[Z_bit] = next_x == 0;
	
	if (((curr_cycle == 1)&(curr_ir == 8'hA8)))
		next_y = curr_a;
	
	if (((curr_cycle == 1)&(curr_ir == 8'hAA)))
		next_x = curr_a;
	
	if (((curr_cycle == 1)&(curr_ir == 8'hB0)))
		next_cycle = (curr_p[C_bit] ? (curr_cycle + 1) : 0);
	
	if (((curr_cycle == 1)&(curr_ir == 8'hB8)))
		next_p[V_bit] = 0;
	
	if (((curr_cycle == 1)&(curr_ir == 8'hBA)))
		next_x = curr_s;
	
	if (((curr_cycle == 2)&(curr_ir == 8'hC4))|
	    ((curr_cycle == 1)&(curr_ir == 8'hC0))|
	    ((curr_cycle == 3)&(curr_ir == 8'hCC)))
		alu_in_lhs = curr_y;
	
	if (((curr_cycle == 2)&((curr_ir == 8'hC5)|(curr_ir == 8'hE4)|(curr_ir == 8'hC4)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hD5)|(curr_ir == 8'hC7)|(curr_ir == 8'hEC)|(curr_ir == 8'hCC)|(curr_ir == 8'hCD)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hD9)|(curr_ir == 8'hD7)|(curr_ir == 8'hDD)|(curr_ir == 8'hCF)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hE0)|(curr_ir == 8'hC0)|(curr_ir == 8'hC9)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hD1)|(curr_ir == 8'hDF)|(curr_ir == 8'hDB)|(curr_ir == 8'hC1)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hD3)|(curr_ir == 8'hC3))))
		next_p[Z_bit] = alu_cmp_z;
	
	if (((curr_cycle == 2)&((curr_ir == 8'hC5)|(curr_ir == 8'hE4)|(curr_ir == 8'hC4)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hD5)|(curr_ir == 8'hC7)|(curr_ir == 8'hEC)|(curr_ir == 8'hCC)|(curr_ir == 8'hCD)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hD9)|(curr_ir == 8'hD7)|(curr_ir == 8'hDD)|(curr_ir == 8'hCF)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hE0)|(curr_ir == 8'hC0)|(curr_ir == 8'hC9)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hD1)|(curr_ir == 8'hDF)|(curr_ir == 8'hDB)|(curr_ir == 8'hC1)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hD3)|(curr_ir == 8'hC3))))
		next_p[N_bit] = alu_cmp_n;
	
	if (((curr_cycle == 2)&((curr_ir == 8'hC5)|(curr_ir == 8'hE4)|(curr_ir == 8'hC4)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hD5)|(curr_ir == 8'hC7)|(curr_ir == 8'hEC)|(curr_ir == 8'hCC)|(curr_ir == 8'hCD)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hD9)|(curr_ir == 8'hD7)|(curr_ir == 8'hDD)|(curr_ir == 8'hCF)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hE0)|(curr_ir == 8'hC0)|(curr_ir == 8'hC9)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hD1)|(curr_ir == 8'hDF)|(curr_ir == 8'hDB)|(curr_ir == 8'hC1)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hD3)|(curr_ir == 8'hC3))))
		next_p[C_bit] = alu_cmp_c;
	
	if (((curr_cycle == 3)&((curr_ir == 8'hD7)|(curr_ir == 8'hCF)))|
	    ((curr_cycle == 2)&(curr_ir == 8'hC7))|
	    ((curr_cycle == 5)&((curr_ir == 8'hC3)|(curr_ir == 8'hD3)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hDF)|(curr_ir == 8'hDB))))
		alu_in_rhs = G_rd_data - 1;
	
	if (((curr_cycle == 5)&((curr_ir == 8'hF7)|(curr_ir == 8'hD7)|(curr_ir == 8'hEF)|(curr_ir == 8'hDF)|(curr_ir == 8'hDB)|(curr_ir == 8'hCF)|(curr_ir == 8'hFF)|(curr_ir == 8'hFB)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hDB)|(curr_ir == 8'hFF)|(curr_ir == 8'hFB)|(curr_ir == 8'hF3)|(curr_ir == 8'hE3)|(curr_ir == 8'hD3)|(curr_ir == 8'hDF)|(curr_ir == 8'hC3)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hE7)|(curr_ir == 8'hD7)|(curr_ir == 8'hF7)|(curr_ir == 8'hEF)|(curr_ir == 8'hC7)|(curr_ir == 8'hCF)))|
	    ((curr_cycle == 7)&((curr_ir == 8'hF3)|(curr_ir == 8'hE3)|(curr_ir == 8'hD3)|(curr_ir == 8'hC3)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hC7)|(curr_ir == 8'hE7))))
		G_wr_data = alu_out_rhs;
	
	if (((curr_cycle == 3)&((curr_ir == 8'hCE)|(curr_ir == 8'hD6)))|
	    ((curr_cycle == 4)&(curr_ir == 8'hDE))|
	    ((curr_cycle == 2)&(curr_ir == 8'hC6)))
		alu_in_rhs = 8'hFF;
	
	if (((curr_cycle == 5)&((curr_ir == 8'hDE)|(curr_ir == 8'hFE)|(curr_ir == 8'hEE)|(curr_ir == 8'hD6)|(curr_ir == 8'hF6)|(curr_ir == 8'hCE)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hF6)|(curr_ir == 8'hCE)|(curr_ir == 8'hD6)|(curr_ir == 8'hEE)|(curr_ir == 8'hC6)|(curr_ir == 8'hE6)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hDE)|(curr_ir == 8'hFE)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hC6)|(curr_ir == 8'hE6))))
		G_wr_data = alu_adc[7:0];
	
	if (((curr_cycle == 6)&((curr_ir == 8'hDE)|(curr_ir == 8'hFE)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hEE)|(curr_ir == 8'hD6)|(curr_ir == 8'hF6)|(curr_ir == 8'hCE)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hC6)|(curr_ir == 8'hE6))))
		next_p[Z_bit] = alu_adc[7:0] == 0;
	
	if (((curr_cycle == 6)&((curr_ir == 8'hDE)|(curr_ir == 8'hFE)))|
	    ((curr_cycle == 5)&((curr_ir == 8'hEE)|(curr_ir == 8'hD6)|(curr_ir == 8'hF6)|(curr_ir == 8'hCE)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hC6)|(curr_ir == 8'hE6))))
		next_p[N_bit] = alu_adc[7];
	
	if (((curr_cycle == 1)&(curr_ir == 8'hC8)))
		next_y = curr_y + 1;
	
	if (((curr_cycle == 1)&(curr_ir == 8'hCA)))
		next_x = curr_x - 1;
	
	if (((curr_cycle == 1)&(curr_ir == 8'hD0)))
		next_cycle = (curr_p[Z_bit] ? 0 : (curr_cycle + 1));
	
	if (((curr_cycle == 1)&(curr_ir == 8'hD8)))
		next_p[D_bit] = 0;
	
	if (((curr_cycle == 2)&(curr_ir == 8'hE4))|
	    ((curr_cycle == 3)&(curr_ir == 8'hEC))|
	    ((curr_cycle == 1)&(curr_ir == 8'hE0)))
		alu_in_lhs = curr_x;
	
	if (((curr_cycle == 5)&((curr_ir == 8'hF1)|(curr_ir == 8'hEF)|(curr_ir == 8'hE1)|(curr_ir == 8'hF7)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hED)|(curr_ir == 8'hF5)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hEB)|(curr_ir == 8'hE9)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hFD)|(curr_ir == 8'hE7)|(curr_ir == 8'hF9)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hFB)|(curr_ir == 8'hFF)))|
	    ((curr_cycle == 7)&((curr_ir == 8'hE3)|(curr_ir == 8'hF3)))|
	    ((curr_cycle == 2)&(curr_ir == 8'hE5)))
		next_a = alu_sbc[7:0];
	
	if (((curr_cycle == 5)&((curr_ir == 8'hF1)|(curr_ir == 8'hEF)|(curr_ir == 8'hE1)|(curr_ir == 8'hF7)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hED)|(curr_ir == 8'hF5)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hEB)|(curr_ir == 8'hE9)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hFD)|(curr_ir == 8'hE7)|(curr_ir == 8'hF9)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hFB)|(curr_ir == 8'hFF)))|
	    ((curr_cycle == 7)&((curr_ir == 8'hE3)|(curr_ir == 8'hF3)))|
	    ((curr_cycle == 2)&(curr_ir == 8'hE5)))
		next_p[C_bit] = alu_sbc_c;
	
	if (((curr_cycle == 5)&((curr_ir == 8'hF1)|(curr_ir == 8'hEF)|(curr_ir == 8'hE1)|(curr_ir == 8'hF7)))|
	    ((curr_cycle == 3)&((curr_ir == 8'hED)|(curr_ir == 8'hF5)))|
	    ((curr_cycle == 1)&((curr_ir == 8'hEB)|(curr_ir == 8'hE9)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hFD)|(curr_ir == 8'hE7)|(curr_ir == 8'hF9)))|
	    ((curr_cycle == 6)&((curr_ir == 8'hFB)|(curr_ir == 8'hFF)))|
	    ((curr_cycle == 7)&((curr_ir == 8'hE3)|(curr_ir == 8'hF3)))|
	    ((curr_cycle == 2)&(curr_ir == 8'hE5)))
		next_p[V_bit] = alu_sbc_v;
	
	if (((curr_cycle == 3)&((curr_ir == 8'hF7)|(curr_ir == 8'hEF)))|
	    ((curr_cycle == 4)&((curr_ir == 8'hFB)|(curr_ir == 8'hFF)))|
	    ((curr_cycle == 2)&(curr_ir == 8'hE7))|
	    ((curr_cycle == 5)&((curr_ir == 8'hF3)|(curr_ir == 8'hE3))))
		alu_in_rhs = G_rd_data + 1;
	
	if (((curr_cycle == 4)&(curr_ir == 8'hFE))|
	    ((curr_cycle == 3)&((curr_ir == 8'hEE)|(curr_ir == 8'hF6)))|
	    ((curr_cycle == 2)&(curr_ir == 8'hE6)))
		alu_in_rhs = 8'h01;
	
	if (((curr_cycle == 1)&(curr_ir == 8'hE8)))
		next_x = curr_x + 1;
	
	if (((curr_cycle == 1)&(curr_ir == 8'hF0)))
		next_cycle = (curr_p[Z_bit] ? (curr_cycle + 1) : 0);
	
	if (((curr_cycle == 1)&(curr_ir == 8'hF8)))
		next_p[D_bit] = 1;
	
	if (((curr_cycle == 0)))
		{next_pch, next_pcl} = force_brk ? curr_pc : curr_pc + 1;
	
	if (((curr_cycle == 0)))
		next_ir = force_brk ? 8'h00 : G_rd_data;
	