
module balloon_fight (I_clock, I_reset, I_phy2, I_prg_addr, I_prg_wren, I_prg_data, O_prg_data, I_chr_addr, I_chr_wren, I_chr_data, O_chr_data, O_ciram_ce, O_ciram_a10, O_ciram_a11, O_irq);
	
	input    wire         I_clock     ;
	input    wire         I_reset     ;
	input    wire         I_phy2      ;
	input    wire[15:0]   I_prg_addr  ;
	input    wire         I_prg_wren  ;
	input    wire[7:0]    I_prg_data  ;
	output   logic[7:0]   O_prg_data  ;
	input    wire[13:0]   I_chr_addr  ;
	input    wire         I_chr_wren  ;
	input    wire[7:0]    I_chr_data  ;
	output   logic[7:0]   O_chr_data  ;
	output   logic        O_ciram_ce  ;
	output   logic        O_ciram_a10 ;
	output   logic        O_ciram_a11 ;
	output   logic        O_irq       ;
	
	bit[7:0] prg_bits [0:16383];
	
	bit[7:0] chr_bits [0:8191];
	
	initial begin
		prg_bits = '{
			8'hA9, 8'h00, 8'h8D, 8'h00, 8'h20, 8'h8D, 8'h01, 8'h20, 8'hAD, 8'h02, 8'h20, 8'h10, 8'hFB, 8'hAD, 8'h02, 8'h20,
			8'h30, 8'hFB, 8'hAD, 8'h02, 8'h20, 8'h10, 8'hFB, 8'h78, 8'hD8, 8'hA2, 8'hFF, 8'h9A, 8'hA2, 8'h12, 8'hA9, 8'h00,
			8'h95, 8'h00, 8'hE8, 8'hD0, 8'hFB, 8'hA2, 8'h02, 8'hBD, 8'hFA, 8'h07, 8'hDD, 8'h82, 8'hC0, 8'hD0, 8'h05, 8'hCA,
			8'h10, 8'hF5, 8'h30, 8'h43, 8'hA2, 8'h00, 8'h8A, 8'h95, 8'h00, 8'h9D, 8'h00, 8'h07, 8'hE8, 8'hD0, 8'hF8, 8'hA9,
			8'h32, 8'h85, 8'h15, 8'hA9, 8'h32, 8'h20, 8'hDE, 8'hD6, 8'hA9, 8'h00, 8'h85, 8'h46, 8'h20, 8'h79, 8'hC5, 8'hC6,
			8'h15, 8'hD0, 8'hF0, 8'hA2, 8'h0E, 8'hBD, 8'h85, 8'hC0, 8'h9D, 8'h29, 8'h06, 8'hCA, 8'h10, 8'hF7, 8'hA2, 8'h04,
			8'hA9, 8'h00, 8'h95, 8'h03, 8'hCA, 8'h10, 8'hF9, 8'hA9, 8'h00, 8'h20, 8'hDE, 8'hD6, 8'hA2, 8'h02, 8'hBD, 8'h82,
			8'hC0, 8'h9D, 8'hFA, 8'h07, 8'hCA, 8'h10, 8'hF7, 8'hA9, 8'h1E, 8'h85, 8'h01, 8'hA9, 8'h90, 8'h85, 8'h00, 8'h4C,
			8'hD4, 8'hF1, 8'h48, 8'h41, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00,
			8'h00, 8'h05, 8'h02, 8'h00, 8'h48, 8'h8A, 8'h48, 8'h98, 8'h48, 8'hA9, 8'h00, 8'h8D, 8'h03, 8'h20, 8'hA9, 8'h02,
			8'h8D, 8'h14, 8'h40, 8'hA5, 8'h52, 8'hC5, 8'h53, 8'hF0, 8'h03, 8'h20, 8'h7C, 8'hC1, 8'h20, 8'h0D, 8'hD6, 8'h20,
			8'h98, 8'hD7, 8'hE6, 8'h19, 8'hA9, 8'h20, 8'h8D, 8'h06, 8'h20, 8'hA9, 8'h00, 8'h8D, 8'h06, 8'h20, 8'hA9, 8'h00,
			8'h8D, 8'h05, 8'h20, 8'h8D, 8'h05, 8'h20, 8'h20, 8'hF7, 8'hFF, 8'hA9, 8'h01, 8'h85, 8'h02, 8'hA5, 8'h16, 8'hF0,
			8'h20, 8'hAD, 8'h02, 8'h20, 8'h30, 8'hFB, 8'hA2, 8'h04, 8'hA0, 8'hC6, 8'h88, 8'hD0, 8'hFD, 8'hCA, 8'hD0, 8'hFA,
			8'hA5, 8'h18, 8'h05, 8'h00, 8'h8D, 8'h00, 8'h20, 8'hA5, 8'h17, 8'h8D, 8'h05, 8'h20, 8'hA9, 8'h00, 8'h8D, 8'h05,
			8'h20, 8'h68, 8'hA8, 8'h68, 8'hAA, 8'h68, 8'h40, 8'h4C, 8'hF7, 8'hC0, 8'hA5, 8'h00, 8'h29, 8'h7F, 8'h8D, 8'h00,
			8'h20, 8'h85, 8'h00, 8'h60, 8'hA5, 8'h00, 8'h09, 8'h80, 8'hD0, 8'hF4, 8'hA9, 8'h00, 8'h48, 8'h20, 8'h65, 8'hF4,
			8'h68, 8'h8D, 8'h01, 8'h20, 8'h60, 8'hA5, 8'h01, 8'hD0, 8'hF3, 8'h20, 8'h54, 8'hC1, 8'hA0, 8'h00, 8'hB9, 8'h57,
			8'h00, 8'h9D, 8'h00, 8'h03, 8'hE8, 8'hC8, 8'hC4, 8'h56, 8'hD0, 8'hF4, 8'h86, 8'h53, 8'h60, 8'hA9, 8'h57, 8'hA0,
			8'h00, 8'h85, 8'h21, 8'h84, 8'h22, 8'h8A, 8'h48, 8'hA0, 8'h02, 8'hB1, 8'h21, 8'h18, 8'h69, 8'h03, 8'h85, 8'h12,
			8'hA6, 8'h53, 8'hA0, 8'h00, 8'hB1, 8'h21, 8'h9D, 8'h00, 8'h03, 8'hE8, 8'hC8, 8'hC4, 8'h12, 8'hD0, 8'hF5, 8'h86,
			8'h53, 8'h68, 8'hAA, 8'h60, 8'hA6, 8'h53, 8'hA9, 8'h00, 8'h85, 8'h12, 8'hA5, 8'h55, 8'h0A, 8'h0A, 8'h0A, 8'h0A,
			8'h26, 8'h12, 8'h0A, 8'h26, 8'h12, 8'h05, 8'h54, 8'h48, 8'hA5, 8'h12, 8'h09, 8'h20, 8'h9D, 8'h00, 8'h03, 8'hE8,
			8'h68, 8'h9D, 8'h00, 8'h03, 8'hE8, 8'hA5, 8'h56, 8'h9D, 8'h00, 8'h03, 8'hE8, 8'h60, 8'h98, 8'h48, 8'h8A, 8'h48,
			8'h20, 8'h88, 8'hC1, 8'h68, 8'hAA, 8'h68, 8'hA8, 8'h60, 8'hA6, 8'h52, 8'hBD, 8'h00, 8'h03, 8'hE8, 8'h85, 8'h50,
			8'h8D, 8'h06, 8'h20, 8'hBD, 8'h00, 8'h03, 8'hE8, 8'h8D, 8'h06, 8'h20, 8'hBC, 8'h00, 8'h03, 8'hE8, 8'hBD, 8'h00,
			8'h03, 8'hE8, 8'h8D, 8'h07, 8'h20, 8'h88, 8'hD0, 8'hF6, 8'hA5, 8'h50, 8'hC9, 8'h3F, 8'hD0, 8'h10, 8'hA9, 8'h3F,
			8'h8D, 8'h06, 8'h20, 8'hA9, 8'h00, 8'h8D, 8'h06, 8'h20, 8'h8D, 8'h06, 8'h20, 8'h8D, 8'h06, 8'h20, 8'h86, 8'h52,
			8'hE4, 8'h53, 8'hD0, 8'hC4, 8'h60, 8'hA9, 8'h20, 8'h85, 8'hF2, 8'h20, 8'h27, 8'hC5, 8'h20, 8'h39, 8'hC5, 8'hA9,
			8'hFF, 8'h85, 8'hCD, 8'hA9, 8'hAD, 8'h85, 8'h23, 8'hA9, 8'hC4, 8'h85, 8'h24, 8'hA9, 8'h80, 8'h85, 8'h91, 8'h8D,
			8'h88, 8'h04, 8'hA9, 8'h70, 8'h85, 8'h9A, 8'h20, 8'h4A, 8'hCD, 8'hA9, 8'h00, 8'h85, 8'h41, 8'h85, 8'hC9, 8'h85,
			8'hCA, 8'h85, 8'hBA, 8'h85, 8'hC5, 8'h85, 8'hC8, 8'h20, 8'hA5, 8'hF4, 8'hA2, 8'h13, 8'hA9, 8'hFF, 8'h9D, 8'h30,
			8'h05, 8'hA9, 8'hF0, 8'h9D, 8'hA4, 8'h04, 8'hCA, 8'h10, 8'hF3, 8'h20, 8'h70, 8'hF4, 8'h20, 8'h91, 8'hE6, 8'hA5,
			8'hC5, 8'hD0, 8'h03, 8'h20, 8'hF9, 8'hC6, 8'hA5, 8'h19, 8'h4A, 8'hB0, 8'h03, 8'h4C, 8'hD0, 8'hC2, 8'hA5, 8'hC5,
			8'hF0, 8'h05, 8'hC6, 8'hC5, 8'h4C, 8'hD0, 8'hC2, 8'hA5, 8'h17, 8'hD0, 8'h06, 8'hA5, 8'h18, 8'h49, 8'h01, 8'h85,
			8'h18, 8'hC6, 8'h17, 8'hAD, 8'h88, 8'h04, 8'hF0, 8'h15, 8'hEE, 8'h88, 8'h04, 8'hAD, 8'h88, 8'h04, 8'hC9, 8'hF0,
			8'h90, 8'h05, 8'hA9, 8'h00, 8'h8D, 8'h88, 8'h04, 8'hA5, 8'hBD, 8'hF0, 8'h02, 8'hE6, 8'h91, 8'hA2, 8'h07, 8'hBD,
			8'h5D, 8'h05, 8'h30, 8'h19, 8'hFE, 8'h67, 8'h05, 8'hBD, 8'h67, 8'h05, 8'hC9, 8'hF8, 8'hD0, 8'h0F, 8'hA9, 8'hFF,
			8'h9D, 8'h5D, 8'h05, 8'hA9, 8'hF0, 8'h9D, 8'h7B, 8'h05, 8'hA9, 8'h00, 8'h8D, 8'hCE, 8'h05, 8'hCA, 8'h10, 8'hDF,
			8'hA2, 8'h13, 8'hBD, 8'h30, 8'h05, 8'h30, 8'h12, 8'hFE, 8'h90, 8'h04, 8'hBD, 8'h90, 8'h04, 8'hC9, 8'hF8, 8'h90,
			8'h08, 8'hA9, 8'hF0, 8'h9D, 8'hA4, 8'h04, 8'h9D, 8'h30, 8'h05, 8'hCA, 8'h10, 8'hE6, 8'hA5, 8'h17, 8'h29, 8'h07,
			8'hD0, 8'h3E, 8'hA6, 8'h88, 8'hCA, 8'h30, 8'h39, 8'hA9, 8'h00, 8'h85, 8'h3E, 8'hA9, 8'h01, 8'h20, 8'hDE, 8'hD6,
			8'hE6, 8'hC9, 8'hA5, 8'hC9, 8'h29, 8'h1F, 8'hD0, 8'h14, 8'hE6, 8'hCA, 8'hA5, 8'hCA, 8'hC9, 8'h0A, 8'hD0, 8'h0C,
			8'hA9, 8'h02, 8'h85, 8'hCA, 8'hA4, 8'hBA, 8'hC8, 8'h98, 8'h29, 8'h03, 8'h85, 8'hBA, 8'hA6, 8'hCA, 8'hBD, 8'hBF,
			8'hC3, 8'h0A, 8'hA8, 8'hB9, 8'hB5, 8'hC3, 8'h85, 8'h25, 8'hB9, 8'hB6, 8'hC3, 8'h85, 8'h26, 8'h20, 8'hB2, 8'hC3,
			8'hA2, 8'h07, 8'hBD, 8'h5D, 8'h05, 8'h30, 8'h18, 8'h20, 8'hCE, 8'hCE, 8'hAD, 8'hCD, 8'h05, 8'hF0, 8'h10, 8'hCE,
			8'hCD, 8'h05, 8'hEE, 8'hCE, 8'h05, 8'h8A, 8'h48, 8'hAD, 8'h59, 8'h05, 8'h20, 8'hDE, 8'hD6, 8'h68, 8'hAA, 8'h20,
			8'h2F, 8'hCE, 8'hCA, 8'h10, 8'hDD, 8'hA2, 8'h13, 8'hBD, 8'h30, 8'h05, 8'h30, 8'h1B, 8'hA5, 8'hC5, 8'hD0, 8'h14,
			8'h20, 8'hB6, 8'hC9, 8'hBD, 8'hA4, 8'h04, 8'hC9, 8'h02, 8'hB0, 8'h03, 8'h20, 8'h4F, 8'hCA, 8'hC9, 8'hD8, 8'h90,
			8'h03, 8'h20, 8'h4F, 8'hCA, 8'h20, 8'h1C, 8'hCB, 8'hA5, 8'h19, 8'h29, 8'h07, 8'h4A, 8'hA8, 8'hB9, 8'hDD, 8'hC9,
			8'h48, 8'hA5, 8'h19, 8'h4A, 8'h8A, 8'h90, 8'h06, 8'h85, 8'h12, 8'hA9, 8'h13, 8'hE5, 8'h12, 8'h0A, 8'h0A, 8'hA8,
			8'h68, 8'h99, 8'hB1, 8'h02, 8'hBD, 8'hA4, 8'h04, 8'h99, 8'hB0, 8'h02, 8'hBD, 8'h90, 8'h04, 8'h99, 8'hB3, 8'h02,
			8'hA9, 8'h00, 8'h99, 8'hB2, 8'h02, 8'hCA, 8'h10, 8'hAF, 8'hAD, 8'hCE, 8'h05, 8'hC9, 8'h14, 8'h90, 8'h20, 8'hE6,
			8'h47, 8'hA9, 8'h00, 8'h20, 8'hDE, 8'hD6, 8'hC6, 8'h47, 8'hA9, 8'h10, 8'h85, 8'hF2, 8'hE6, 8'hC8, 8'h20, 8'hED,
			8'hD3, 8'h20, 8'h27, 8'hC5, 8'hC6, 8'hC8, 8'hA2, 8'h64, 8'h20, 8'h5E, 8'hF4, 8'hA9, 8'h20, 8'h85, 8'hF2, 8'hA2,
			8'hF0, 8'hAD, 8'h88, 8'h04, 8'hF0, 8'h02, 8'hA2, 8'h88, 8'h8E, 8'h00, 8'h02, 8'h8E, 8'h04, 8'h02, 8'h8D, 8'h03,
			8'h02, 8'h18, 8'h69, 8'h08, 8'h8D, 8'h07, 8'h02, 8'hA5, 8'h19, 8'h29, 8'h03, 8'h8D, 8'h02, 8'h02, 8'h8D, 8'h06,
			8'h02, 8'hA2, 8'hE3, 8'h8E, 8'h01, 8'h02, 8'hE8, 8'h8E, 8'h05, 8'h02, 8'hA5, 8'h88, 8'h30, 8'h03, 8'h4C, 8'h09,
			8'hC2, 8'h20, 8'h79, 8'hC5, 8'hA9, 8'h01, 8'h85, 8'hF0, 8'h20, 8'h65, 8'hF4, 8'hA9, 8'h02, 8'h85, 8'hF2, 8'h4C,
			8'h6A, 8'hF3, 8'h6C, 8'h25, 8'h00, 8'hC9, 8'hC3, 8'hF7, 8'hC3, 8'h3E, 8'hC4, 8'h5F, 8'hC4, 8'h5E, 8'hC4, 8'h00,
			8'h00, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h04, 8'h03, 8'h01, 8'hA0, 8'h00, 8'hB1, 8'h23, 8'hE6, 8'h23, 8'hD0,
			8'h02, 8'hE6, 8'h24, 8'hAA, 8'hF0, 8'h20, 8'h0A, 8'h0A, 8'h0A, 8'h85, 8'h15, 8'hA9, 8'h00, 8'h85, 8'h14, 8'h8A,
			8'h29, 8'hC0, 8'hC9, 8'h80, 8'hD0, 8'h06, 8'h20, 8'h6B, 8'hC4, 8'h4C, 8'hC9, 8'hC3, 8'hC9, 8'h00, 8'hD0, 8'h06,
			8'h20, 8'h86, 8'hC4, 8'h4C, 8'hC9, 8'hC3, 8'h60, 8'h20, 8'hB3, 8'hF1, 8'h29, 8'h7F, 8'hC9, 8'h04, 8'h90, 8'h0C,
			8'hC9, 8'h18, 8'hB0, 8'h08, 8'h0A, 8'h0A, 8'h0A, 8'h85, 8'h15, 8'h20, 8'h6B, 8'hC4, 8'h20, 8'hB3, 8'hF1, 8'h29,
			8'h3F, 8'hC9, 8'h02, 8'h90, 8'h24, 8'hC9, 8'h18, 8'hB0, 8'h20, 8'h0A, 8'h0A, 8'h0A, 8'h85, 8'h15, 8'h20, 8'hB3,
			8'hF1, 8'h29, 8'h3F, 8'hA6, 8'hBA, 8'h7D, 8'h3A, 8'hC4, 8'h85, 8'h14, 8'h20, 8'h86, 8'hC4, 8'h20, 8'hB3, 8'hF1,
			8'h4A, 8'h90, 8'hD9, 8'h20, 8'h4F, 8'hCA, 8'h4C, 8'h0C, 8'hC4, 8'h60, 8'h20, 8'h30, 8'h40, 8'h60, 8'h20, 8'hB3,
			8'hF1, 8'h29, 8'hCF, 8'hD0, 8'hB2, 8'hA4, 8'h89, 8'hC8, 8'hD0, 8'hAD, 8'hA9, 8'hE6, 8'h85, 8'h9B, 8'hA5, 8'h1B,
			8'h29, 8'h7F, 8'h69, 8'h40, 8'h85, 8'h92, 8'hA9, 8'h80, 8'h85, 8'h89, 8'hA9, 8'h00, 8'h85, 8'h80, 8'h60, 8'h20,
			8'h0C, 8'hC4, 8'h20, 8'hB3, 8'hF1, 8'h29, 8'h7F, 8'h9D, 8'h08, 8'h05, 8'h60, 8'hA2, 8'h07, 8'hBD, 8'h5D, 8'h05,
			8'h30, 8'h04, 8'hCA, 8'h10, 8'hF8, 8'h60, 8'hA9, 8'h01, 8'h9D, 8'h5D, 8'h05, 8'hA9, 8'h00, 8'h9D, 8'h67, 8'h05,
			8'hA5, 8'h15, 8'h9D, 8'h7B, 8'h05, 8'h60, 8'hA2, 8'h13, 8'hBD, 8'h30, 8'h05, 8'h30, 8'h04, 8'hCA, 8'h10, 8'hF8,
			8'h60, 8'hA9, 8'h00, 8'h9D, 8'h30, 8'h05, 8'h9D, 8'h90, 8'h04, 8'h9D, 8'hF4, 8'h04, 8'h9D, 8'h08, 8'h05, 8'h9D,
			8'hE0, 8'h04, 8'hA5, 8'h14, 8'h9D, 8'h1C, 8'h05, 8'hA5, 8'h15, 8'h9D, 8'hA4, 8'h04, 8'h60, 8'h00, 8'h00, 8'h09,
			8'h00, 8'h08, 8'h8C, 8'h00, 8'h07, 8'h18, 8'h00, 8'h18, 8'h00, 8'h19, 8'h00, 8'h1A, 8'h00, 8'h84, 8'h94, 8'h1A,
			8'h00, 8'h1A, 8'h00, 8'h1A, 8'h00, 8'h0B, 8'h12, 8'h00, 8'h0C, 8'h13, 8'h00, 8'h0D, 8'h14, 8'h00, 8'h14, 8'h00,
			8'h00, 8'h90, 8'h00, 8'h07, 8'h00, 8'h07, 8'h8C, 8'h96, 8'h00, 8'h08, 8'h00, 8'h09, 8'h00, 8'h00, 8'h18, 8'h00,
			8'h17, 8'h00, 8'h16, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h8A, 8'h90, 8'h00, 8'h00, 8'h00, 8'h08, 8'h00,
			8'h09, 8'h98, 8'h00, 8'h0A, 8'h00, 8'h00, 8'h00, 8'h86, 8'h8A, 8'h15, 8'h00, 8'h14, 8'h00, 8'h8E, 8'h13, 8'h00,
			8'h00, 8'h03, 8'h0D, 8'h00, 8'h0D, 8'h0E, 8'h00, 8'h0C, 8'h0D, 8'h00, 8'h0D, 8'h19, 8'h00, 8'h86, 8'h92, 8'h00,
			8'h00, 8'h98, 8'h00, 8'h00, 8'h0A, 8'h12, 8'h00, 8'h09, 8'h13, 8'h00, 8'h08, 8'h14, 8'h00, 8'h07, 8'h15, 8'h00,
			8'h07, 8'h16, 8'h00, 8'h07, 8'h00, 8'h00, 8'h00, 8'h20, 8'hE2, 8'hD0, 8'h0E, 8'h59, 8'h05, 8'hAD, 8'h59, 8'h05,
			8'h0A, 8'h0A, 8'h6D, 8'h59, 8'h05, 8'h8D, 8'h59, 8'h05, 8'h60, 8'hA9, 8'h00, 8'h85, 8'h12, 8'hA5, 8'h12, 8'h0A,
			8'h0A, 8'h65, 8'h12, 8'h85, 8'h1D, 8'hA9, 8'h07, 8'h85, 8'h1E, 8'hA0, 8'h04, 8'hB1, 8'h1D, 8'hD9, 8'h03, 8'h00,
			8'h90, 8'h11, 8'hD0, 8'h05, 8'h88, 8'h10, 8'hF4, 8'h30, 8'h0A, 8'hE6, 8'h12, 8'hA5, 8'h12, 8'hC9, 8'h32, 8'hD0,
			8'hDC, 8'hC6, 8'h12, 8'hE6, 8'h12, 8'hA5, 8'h12, 8'h48, 8'h85, 8'h43, 8'hA0, 8'h0A, 8'h20, 8'h7C, 8'hD7, 8'h85,
			8'h4A, 8'hA5, 8'h43, 8'h85, 8'h49, 8'h68, 8'h85, 8'h12, 8'h60, 8'h20, 8'h39, 8'hC5, 8'hC6, 8'h12, 8'hA9, 8'h31,
			8'h38, 8'hE5, 8'h12, 8'h85, 8'h13, 8'h0A, 8'h0A, 8'h65, 8'h13, 8'hA8, 8'hA5, 8'h12, 8'h0A, 8'h0A, 8'h65, 8'h12,
			8'h85, 8'h1D, 8'h18, 8'h69, 8'h05, 8'h85, 8'h1F, 8'hA9, 8'h07, 8'h85, 8'h1E, 8'h85, 8'h20, 8'h98, 8'hF0, 8'h0C,
			8'h88, 8'hB1, 8'h1D, 8'h91, 8'h1F, 8'h88, 8'hD0, 8'hF9, 8'hB1, 8'h1D, 8'h91, 8'h1F, 8'hA0, 8'h04, 8'hB9, 8'h03,
			8'h00, 8'h91, 8'h1D, 8'h88, 8'h10, 8'hF8, 8'h60, 8'h01, 8'h02, 8'h03, 8'h03, 8'h02, 8'h01, 8'hFF, 8'h03, 8'h04,
			8'h05, 8'h06, 8'hFF, 8'hAD, 8'h8D, 8'h04, 8'h4A, 8'h4A, 8'h4A, 8'hAA, 8'hAD, 8'h8A, 8'h04, 8'hD0, 8'h06, 8'hBD,
			8'hB7, 8'hC5, 8'h4C, 8'hD8, 8'hC5, 8'hBD, 8'hBB, 8'hC5, 8'h85, 8'h87, 8'hA2, 8'h08, 8'h20, 8'hA4, 8'hE3, 8'hAD,
			8'h8C, 8'h04, 8'hF0, 8'h2F, 8'hAE, 8'h8B, 8'h04, 8'hAD, 8'h8D, 8'h04, 8'hC9, 8'h20, 8'hD0, 8'h06, 8'hA9, 8'hFF,
			8'h95, 8'h88, 8'h30, 8'h1C, 8'hB0, 8'h1D, 8'hAD, 8'h50, 8'h04, 8'hD0, 8'h07, 8'hA5, 8'h99, 8'h18, 8'h69, 8'h04,
			8'hD0, 8'h05, 8'hA5, 8'h99, 8'h38, 8'hE9, 8'h04, 8'h95, 8'h91, 8'hA5, 8'hA2, 8'h38, 8'hE9, 8'h0A, 8'h95, 8'h9A,
			8'h20, 8'hA4, 8'hE3, 8'h60, 8'hA9, 8'hFF, 8'h8D, 8'h8B, 8'h04, 8'hA2, 8'h07, 8'hB5, 8'h88, 8'h30, 8'h0C, 8'hB5,
			8'h9A, 8'hC9, 8'hB4, 8'h90, 8'h06, 8'hB5, 8'h91, 8'hC5, 8'h99, 8'hF0, 8'h04, 8'hCA, 8'h10, 8'hED, 8'h60, 8'h8E,
			8'h8B, 8'h04, 8'hBD, 8'h48, 8'h04, 8'h8D, 8'h50, 8'h04, 8'hA9, 8'h00, 8'h8D, 8'h8A, 8'h04, 8'h8D, 8'h8D, 8'h04,
			8'h8D, 8'h8C, 8'h04, 8'h8D, 8'h89, 8'h04, 8'hA9, 8'hDC, 8'h85, 8'hA2, 8'h60, 8'hE6, 8'h99, 8'hA5, 8'h99, 8'hC9,
			8'hB1, 8'h90, 8'h04, 8'hA9, 8'h40, 8'h85, 8'h99, 8'h60, 8'hAD, 8'h89, 8'h04, 8'hD0, 8'h12, 8'hC6, 8'hA2, 8'hA5,
			8'hA2, 8'hC9, 8'hC4, 8'hB0, 8'h0C, 8'hE6, 8'hA2, 8'hEE, 8'h8A, 8'h04, 8'hEE, 8'h89, 8'h04, 8'hD0, 8'h02, 8'hE6,
			8'hA2, 8'hEE, 8'h8D, 8'h04, 8'hAD, 8'h8D, 8'h04, 8'hC9, 8'h18, 8'hD0, 8'h28, 8'hAE, 8'h8B, 8'h04, 8'hB5, 8'h88,
			8'h30, 8'h21, 8'hB5, 8'h9A, 8'h18, 8'h69, 8'h10, 8'hC5, 8'hA2, 8'h90, 8'h18, 8'hBC, 8'h51, 8'h04, 8'hB9, 8'hB8,
			8'hC6, 8'h9D, 8'h51, 8'h04, 8'hA9, 8'h00, 8'h95, 8'h7F, 8'h95, 8'h88, 8'hA5, 8'hF2, 8'h09, 8'h40, 8'h85, 8'hF2,
			8'hEE, 8'h8C, 8'h04, 8'hAD, 8'h8A, 8'h04, 8'hF0, 8'h0F, 8'hAD, 8'h8D, 8'h04, 8'hC9, 8'h28, 8'hF0, 8'h04, 8'hC9,
			8'h30, 8'hD0, 8'h04, 8'hA9, 8'hCC, 8'h85, 8'hA2, 8'h60, 8'h08, 8'h09, 8'h0A, 8'h0B, 8'h08, 8'h09, 8'h0A, 8'h0B,
			8'h08, 8'h09, 8'h0A, 8'h0B, 8'hAD, 8'h89, 8'h04, 8'hD0, 8'h2F, 8'hAE, 8'h8B, 8'h04, 8'hB5, 8'h88, 8'h30, 8'h10,
			8'hB5, 8'h9A, 8'hC9, 8'hB4, 8'h90, 8'h0A, 8'hB5, 8'h91, 8'hC9, 8'h40, 8'h90, 8'h04, 8'hC9, 8'hB1, 8'h90, 8'h0E,
			8'hA9, 8'h30, 8'h38, 8'hED, 8'h8D, 8'h04, 8'h8D, 8'h8D, 8'h04, 8'hEE, 8'h89, 8'h04, 8'hD0, 8'h0A, 8'hB5, 8'h91,
			8'h85, 8'h99, 8'hBD, 8'h48, 8'h04, 8'h8D, 8'h50, 8'h04, 8'h60, 8'hA5, 8'h87, 8'h10, 8'h10, 8'h20, 8'h4B, 8'hC6,
			8'h20, 8'h14, 8'hC6, 8'hAD, 8'h8B, 8'h04, 8'h10, 8'h01, 8'h60, 8'hA9, 8'h40, 8'h85, 8'hF3, 8'h20, 8'hC4, 8'hC6,
			8'h20, 8'h58, 8'hC6, 8'h4C, 8'hC3, 8'hC5, 8'hA2, 8'h01, 8'hA9, 8'hFF, 8'h9D, 8'h30, 8'h05, 8'h9D, 8'h44, 8'h05,
			8'hCA, 8'h10, 8'hF5, 8'h20, 8'h7A, 8'hC7, 8'hA6, 8'h3C, 8'hE0, 8'h18, 8'h90, 8'h02, 8'hA2, 8'h18, 8'hBD, 8'h48,
			8'hC7, 8'h85, 8'hBA, 8'hBD, 8'h61, 8'hC7, 8'h85, 8'hB8, 8'hA9, 8'hF0, 8'h8D, 8'hE0, 8'h02, 8'h8D, 8'hE4, 8'h02,
			8'h8D, 8'hE8, 8'h02, 8'hA9, 8'h03, 8'h4C, 8'h56, 8'hC8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h02, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01,
			8'h01, 8'h0F, 8'h0F, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0C, 8'h0C, 8'h0A, 8'h0A, 8'h0A,
			8'h08, 8'h0A, 8'h0A, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h05, 8'hA5, 8'hA3, 8'h10, 8'h03, 8'h85, 8'hA4,
			8'h60, 8'h20, 8'hB3, 8'hF1, 8'hC5, 8'hA3, 8'h90, 8'hF6, 8'hF0, 8'hF4, 8'h18, 8'hE5, 8'hA3, 8'h4C, 8'h84, 8'hC7,
			8'hA5, 8'h19, 8'h29, 8'h7F, 8'hF0, 8'h01, 8'h60, 8'hC6, 8'hB8, 8'hD0, 8'hFB, 8'hA2, 8'h00, 8'hBD, 8'h30, 8'h05,
			8'h30, 8'h0B, 8'hE8, 8'hBD, 8'h30, 8'h05, 8'h30, 8'h05, 8'hA9, 8'h01, 8'h85, 8'hB8, 8'h60, 8'hA4, 8'hA4, 8'h84,
			8'hA5, 8'h10, 8'h01, 8'h60, 8'hA9, 8'h80, 8'h9D, 8'hB8, 8'h04, 8'h9D, 8'hCC, 8'h04, 8'hA9, 8'h00, 8'h9D, 8'h30,
			8'h05, 8'hB9, 8'hB2, 8'h00, 8'h9D, 8'h90, 8'h04, 8'hB9, 8'hB5, 8'h00, 8'h9D, 8'hA4, 8'h04, 8'hA4, 8'hBA, 8'h20,
			8'hB3, 8'hF1, 8'h29, 8'h1F, 8'h79, 8'h9F, 8'hC8, 8'h9D, 8'h08, 8'h05, 8'hB9, 8'hAB, 8'hC8, 8'h9D, 8'h1C, 8'h05,
			8'hB9, 8'hA5, 8'hC8, 8'h9D, 8'hE0, 8'h04, 8'hB9, 8'hB1, 8'hC8, 8'h9D, 8'hF4, 8'h04, 8'h20, 8'hB3, 8'hF1, 8'h29,
			8'h03, 8'h9D, 8'h44, 8'h05, 8'hA8, 8'hB9, 8'h97, 8'hC8, 8'h18, 8'h7D, 8'h90, 8'h04, 8'h9D, 8'h90, 8'h04, 8'hB9,
			8'h9B, 8'hC8, 8'h18, 8'h7D, 8'hA4, 8'h04, 8'h9D, 8'hA4, 8'h04, 8'hB9, 8'h8F, 8'hC8, 8'hF0, 8'h03, 8'h20, 8'h3D,
			8'hCA, 8'hB9, 8'h93, 8'hC8, 8'hF0, 8'h03, 8'h20, 8'h55, 8'hCA, 8'hA5, 8'hBA, 8'hC9, 8'h05, 8'hB0, 8'h02, 8'hE6,
			8'hBA, 8'hA9, 8'h06, 8'h38, 8'hE5, 8'hBA, 8'h85, 8'hB8, 8'hA5, 8'hF0, 8'h09, 8'h04, 8'h85, 8'hF0, 8'h4C, 8'h7A,
			8'hC7, 8'hA5, 8'hB8, 8'hC9, 8'h01, 8'hD0, 8'h53, 8'hAD, 8'h30, 8'h05, 8'h30, 8'h0A, 8'hAD, 8'h31, 8'h05, 8'h30,
			8'h05, 8'hA9, 8'h02, 8'h85, 8'hB8, 8'h60, 8'hA5, 8'h19, 8'h29, 8'h7F, 8'hC9, 8'h40, 8'h90, 8'h3C, 8'hD0, 8'h06,
			8'hA5, 8'hF1, 8'h09, 8'h08, 8'h85, 8'hF1, 8'h29, 8'h03, 8'hAA, 8'hBD, 8'h8B, 8'hC8, 8'h85, 8'h5A, 8'hA6, 8'hA4,
			8'h30, 8'h28, 8'hA9, 8'h23, 8'h85, 8'h57, 8'hB5, 8'hA6, 8'h85, 8'h58, 8'hA9, 8'h01, 8'h85, 8'h59, 8'h20, 8'h83,
			8'hC8, 8'hB5, 8'hA9, 8'h85, 8'h58, 8'h20, 8'h83, 8'hC8, 8'hB5, 8'hAC, 8'h85, 8'h58, 8'h20, 8'h83, 8'hC8, 8'hB5,
			8'hAF, 8'h85, 8'h58, 8'hA9, 8'h57, 8'hA0, 8'h00, 8'h4C, 8'h31, 8'hC1, 8'h60, 8'h55, 8'hFF, 8'h00, 8'hFF, 8'h00,
			8'h00, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'h10, 8'h10, 8'hF0, 8'hF0, 8'hDE, 8'h22, 8'h22, 8'hDE, 8'h60,
			8'h70, 8'h80, 8'h90, 8'hA0, 8'hB0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hF0, 8'h20, 8'h50, 8'h80,
			8'hB0, 8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h01, 8'hA2, 8'h01, 8'hBD, 8'h30, 8'h05, 8'h10, 8'h03, 8'h4C, 8'hAF,
			8'hC9, 8'hBD, 8'h44, 8'h05, 8'h30, 8'h7B, 8'hA8, 8'h8A, 8'h48, 8'hA6, 8'hA5, 8'hB5, 8'hB2, 8'h79, 8'hE5, 8'hC9,
			8'h8D, 8'hE3, 8'h02, 8'h8D, 8'hE7, 8'h02, 8'h8D, 8'hEB, 8'h02, 8'hB5, 8'hB5, 8'h79, 8'hF5, 8'hC9, 8'h8D, 8'hE0,
			8'h02, 8'h79, 8'h05, 8'hCA, 8'h8D, 8'hE4, 8'h02, 8'h79, 8'h05, 8'hCA, 8'h8D, 8'hE8, 8'h02, 8'h98, 8'h29, 8'h03,
			8'hAA, 8'h98, 8'h4A, 8'h4A, 8'hA8, 8'hA5, 8'h19, 8'h4A, 8'h4A, 8'hB0, 8'h04, 8'h98, 8'h69, 8'h05, 8'hA8, 8'hB9,
			8'h15, 8'hCA, 8'h8D, 8'hE1, 8'h02, 8'hB9, 8'h1F, 8'hCA, 8'h8D, 8'hE5, 8'h02, 8'hB9, 8'h29, 8'hCA, 8'h8D, 8'hE9,
			8'h02, 8'hBD, 8'h33, 8'hCA, 8'h8D, 8'hE2, 8'h02, 8'h8D, 8'hE6, 8'h02, 8'h8D, 8'hEA, 8'h02, 8'h68, 8'hAA, 8'hA5,
			8'h19, 8'h29, 8'h07, 8'hD0, 8'h12, 8'hBD, 8'h44, 8'h05, 8'h18, 8'h69, 8'h04, 8'h9D, 8'h44, 8'h05, 8'hC9, 8'h14,
			8'h90, 8'h05, 8'hA9, 8'hFF, 8'h9D, 8'h44, 8'h05, 8'hBD, 8'h44, 8'h05, 8'hC9, 8'h10, 8'hB0, 8'h03, 8'h4C, 8'hAF,
			8'hC9, 8'h20, 8'hB6, 8'hC9, 8'hBD, 8'h90, 8'h04, 8'hC9, 8'h02, 8'hB0, 8'h03, 8'h20, 8'h37, 8'hCA, 8'hBD, 8'h90,
			8'h04, 8'hC9, 8'hF7, 8'h90, 8'h03, 8'h20, 8'h37, 8'hCA, 8'hBD, 8'hA4, 8'h04, 8'hC9, 8'h02, 8'hB0, 8'h03, 8'h20,
			8'h4F, 8'hCA, 8'hBD, 8'hA4, 8'h04, 8'hC9, 8'hE0, 8'h90, 8'h0D, 8'hA9, 8'hFF, 8'h9D, 8'h30, 8'h05, 8'hA9, 8'hF0,
			8'h9D, 8'hA4, 8'h04, 8'h4C, 8'hAF, 8'hC9, 8'h20, 8'h67, 8'hCA, 8'h20, 8'h1C, 8'hCB, 8'hBC, 8'h30, 8'h05, 8'hC8,
			8'h98, 8'h29, 8'h07, 8'h9D, 8'h30, 8'h05, 8'hBC, 8'h30, 8'h05, 8'hB9, 8'hDD, 8'hC9, 8'h85, 8'h12, 8'h8A, 8'h0A,
			8'h0A, 8'h18, 8'hA8, 8'hBD, 8'hA4, 8'h04, 8'hC9, 8'hD0, 8'h99, 8'h00, 8'h02, 8'hBD, 8'h90, 8'h04, 8'h99, 8'h03,
			8'h02, 8'hA5, 8'h12, 8'h99, 8'h01, 8'h02, 8'hA9, 8'h00, 8'h90, 8'h02, 8'hA9, 8'h20, 8'h99, 8'h02, 8'h02, 8'hCA,
			8'h30, 8'h03, 8'h4C, 8'hB9, 8'hC8, 8'h60, 8'hBD, 8'h08, 8'h05, 8'h18, 8'h7D, 8'hB8, 8'h04, 8'h9D, 8'hB8, 8'h04,
			8'hBD, 8'hE0, 8'h04, 8'h7D, 8'h90, 8'h04, 8'h9D, 8'h90, 8'h04, 8'hBD, 8'h1C, 8'h05, 8'h18, 8'h7D, 8'hCC, 8'h04,
			8'h9D, 8'hCC, 8'h04, 8'hBD, 8'hF4, 8'h04, 8'h7D, 8'hA4, 8'h04, 8'h9D, 8'hA4, 8'h04, 8'h60, 8'h9D, 8'h9E, 8'h9F,
			8'h9E, 8'h9D, 8'hA0, 8'hA1, 8'hA0, 8'h08, 8'h08, 8'hF0, 8'hF0, 8'h08, 8'h08, 8'hF0, 8'hF0, 8'h08, 8'h08, 8'hF0,
			8'hF0, 8'h08, 8'h08, 8'hF0, 8'hF0, 8'hEE, 8'h0A, 8'h0A, 8'hEE, 8'hEE, 8'h0A, 8'h0A, 8'hEE, 8'hEE, 8'h0A, 8'h0A,
			8'hEE, 8'hEE, 8'h0A, 8'h0A, 8'hEE, 8'hF8, 8'h08, 8'h08, 8'hF8, 8'hF8, 8'h08, 8'h08, 8'hF8, 8'hF8, 8'h08, 8'h08,
			8'hF8, 8'hF8, 8'h08, 8'h08, 8'hF8, 8'h91, 8'h93, 8'h97, 8'h97, 8'hFC, 8'h92, 8'h95, 8'h9A, 8'h9A, 8'hFC, 8'hFC,
			8'h94, 8'h98, 8'h98, 8'hFC, 8'hFC, 8'h96, 8'h9B, 8'h9B, 8'hFC, 8'hFC, 8'hFC, 8'h99, 8'h99, 8'hFC, 8'hFC, 8'hFC,
			8'h9C, 8'h9C, 8'hFC, 8'hC0, 8'h40, 8'h00, 8'h80, 8'hA5, 8'hF3, 8'h09, 8'h80, 8'h85, 8'hF3, 8'hA9, 8'h00, 8'h38,
			8'hFD, 8'h08, 8'h05, 8'h9D, 8'h08, 8'h05, 8'hA9, 8'h00, 8'hFD, 8'hE0, 8'h04, 8'h9D, 8'hE0, 8'h04, 8'h60, 8'hA5,
			8'hF3, 8'h09, 8'h80, 8'h85, 8'hF3, 8'hA9, 8'h00, 8'h38, 8'hFD, 8'h1C, 8'h05, 8'h9D, 8'h1C, 8'h05, 8'hA9, 8'h00,
			8'hFD, 8'hF4, 8'h04, 8'h9D, 8'hF4, 8'h04, 8'h60, 8'hA4, 8'hCD, 8'hA9, 8'h00, 8'h85, 8'hCC, 8'hB1, 8'h27, 8'h38,
			8'hE9, 8'h08, 8'hDD, 8'hA4, 8'h04, 8'hB0, 8'h66, 8'h69, 8'h03, 8'hDD, 8'hA4, 8'h04, 8'h90, 8'h04, 8'hA9, 8'h01,
			8'hD0, 8'h10, 8'hB1, 8'h29, 8'hDD, 8'hA4, 8'h04, 8'h90, 8'h54, 8'hE9, 8'h03, 8'hDD, 8'hA4, 8'h04, 8'hB0, 8'h1D,
			8'hA9, 8'h02, 8'h85, 8'hCC, 8'hB1, 8'h23, 8'hC9, 8'h10, 8'hF0, 8'h08, 8'h38, 8'hE9, 8'h04, 8'hDD, 8'h90, 8'h04,
			8'hB0, 8'h07, 8'hB1, 8'h25, 8'hDD, 8'h90, 8'h04, 8'hB0, 8'h04, 8'hA9, 8'h00, 8'h85, 8'hCC, 8'hB1, 8'h23, 8'hC9,
			8'h10, 8'hF0, 8'h15, 8'h38, 8'hE9, 8'h08, 8'hDD, 8'h90, 8'h04, 8'hB0, 8'h22, 8'h69, 8'h03, 8'hDD, 8'h90, 8'h04,
			8'h90, 8'h06, 8'hA5, 8'hCC, 8'h09, 8'h04, 8'hD0, 8'h13, 8'hB1, 8'h25, 8'hC9, 8'hFF, 8'hF0, 8'h0F, 8'hDD, 8'h90,
			8'h04, 8'h90, 8'h0A, 8'hE9, 8'h03, 8'hB0, 8'h06, 8'hA5, 8'hCC, 8'h09, 8'h08, 8'h85, 8'hCC, 8'hA5, 8'hCC, 8'hD0,
			8'h07, 8'h88, 8'h30, 8'h03, 8'h4C, 8'h69, 8'hCA, 8'h60, 8'h46, 8'hCC, 8'h90, 8'h08, 8'hBD, 8'hF4, 8'h04, 8'h30,
			8'h03, 8'h20, 8'h4F, 8'hCA, 8'h46, 8'hCC, 8'h90, 8'h08, 8'hBD, 8'hF4, 8'h04, 8'h10, 8'h03, 8'h20, 8'h4F, 8'hCA,
			8'h46, 8'hCC, 8'h90, 8'h08, 8'hBD, 8'hE0, 8'h04, 8'h30, 8'h03, 8'h20, 8'h37, 8'hCA, 8'h46, 8'hCC, 8'h90, 8'h08,
			8'hBD, 8'hE0, 8'h04, 8'h10, 8'h03, 8'h20, 8'h37, 8'hCA, 8'h4C, 8'hE1, 8'hCA, 8'h60, 8'hA0, 8'h01, 8'hB9, 8'h88,
			8'h00, 8'h30, 8'h4D, 8'hF0, 8'h4B, 8'hB9, 8'hBD, 8'h00, 8'hD0, 8'h46, 8'hBD, 8'h90, 8'h04, 8'h38, 8'hF9, 8'h91,
			8'h00, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h08, 8'hB0, 8'h38, 8'hBD, 8'hA4, 8'h04, 8'h38, 8'hF9, 8'h9A, 8'h00, 8'h38,
			8'hE9, 8'h08, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h0C, 8'hB0, 8'h27, 8'hA9, 8'h00, 8'h99, 8'h88, 8'h00, 8'hA9, 8'h01,
			8'h99, 8'h7F, 8'h00, 8'h99, 8'hC1, 8'h00, 8'hA9, 8'h0B, 8'h99, 8'h51, 8'h04, 8'hA9, 8'h20, 8'h99, 8'h5A, 8'h04,
			8'hA5, 8'hF0, 8'h09, 8'h80, 8'h85, 8'hF0, 8'hA9, 8'hF0, 8'h9D, 8'hA4, 8'h04, 8'hA9, 8'hFF, 8'h9D, 8'h30, 8'h05,
			8'h88, 8'h10, 8'hAB, 8'h60, 8'hAE, 8'hD1, 8'h05, 8'h30, 8'h2E, 8'h20, 8'hA8, 8'hCB, 8'hBD, 8'h04, 8'h06, 8'hF0,
			8'h23, 8'h8A, 8'h45, 8'h19, 8'h29, 8'h01, 8'hD0, 8'h1C, 8'hBC, 8'hFA, 8'h05, 8'hC8, 8'h98, 8'h29, 8'h03, 8'h9D,
			8'hFA, 8'h05, 8'h20, 8'hCB, 8'hCC, 8'hBD, 8'hFA, 8'h05, 8'hC9, 8'h01, 8'hD0, 8'h08, 8'hDE, 8'h0E, 8'h06, 8'hD0,
			8'h03, 8'hDE, 8'h04, 8'h06, 8'hCA, 8'h10, 8'hD2, 8'h60, 8'hA0, 8'h07, 8'hBD, 8'h04, 8'h06, 8'hD0, 8'h03, 8'h4C,
			8'h3A, 8'hCC, 8'hB9, 8'h88, 8'h00, 8'h30, 8'h78, 8'hF0, 8'h76, 8'hC0, 8'h02, 8'h90, 8'h04, 8'hC9, 8'h01, 8'hF0,
			8'h6E, 8'hB9, 8'h91, 8'h00, 8'h18, 8'h69, 8'h08, 8'h38, 8'hFD, 8'hD2, 8'h05, 8'h85, 8'h12, 8'h20, 8'h8E, 8'hF0,
			8'hC9, 8'h12, 8'hB0, 8'h5B, 8'hB9, 8'h9A, 8'h00, 8'h18, 8'h69, 8'h0C, 8'h38, 8'hFD, 8'hDC, 8'h05, 8'h85, 8'h13,
			8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h12, 8'hB0, 8'h48, 8'hA5, 8'h12, 8'h30, 8'h11, 8'hC9, 8'h03, 8'h90, 8'h1C, 8'hA9,
			8'h02, 8'h99, 8'h1B, 8'h04, 8'h20, 8'h33, 8'hCC, 8'h20, 8'hBB, 8'hEB, 8'hD0, 8'h0F, 8'hC9, 8'hFD, 8'hB0, 8'h0B,
			8'hA9, 8'hFE, 8'h99, 8'h1B, 8'h04, 8'h20, 8'hBB, 8'hEB, 8'h20, 8'h33, 8'hCC, 8'hA5, 8'h13, 8'h30, 8'h11, 8'hC9,
			8'h03, 8'h90, 8'h1C, 8'hA9, 8'h02, 8'h99, 8'h2D, 8'h04, 8'h20, 8'hB2, 8'hEB, 8'h20, 8'h33, 8'hCC, 8'hD0, 8'h0F,
			8'hC9, 8'hFD, 8'hB0, 8'h0B, 8'hA9, 8'hFE, 8'h99, 8'h2D, 8'h04, 8'h20, 8'hB2, 8'hEB, 8'h20, 8'h33, 8'hCC, 8'h88,
			8'h10, 8'h80, 8'h60, 8'hA5, 8'hF1, 8'h09, 8'h02, 8'h85, 8'hF1, 8'h60, 8'hB9, 8'h88, 8'h00, 8'h30, 8'h79, 8'hF0,
			8'h77, 8'hC0, 8'h02, 8'h90, 8'h2E, 8'hBD, 8'hFA, 8'h05, 8'hC9, 8'h03, 8'hD0, 8'h27, 8'hBD, 8'hD2, 8'h05, 8'h38,
			8'hE9, 8'h0A, 8'hD9, 8'h91, 8'h00, 8'hB0, 8'h1C, 8'h69, 8'h04, 8'hD9, 8'h91, 8'h00, 8'h90, 8'h15, 8'hBD, 8'hDC,
			8'h05, 8'h38, 8'hE9, 8'h1C, 8'hD9, 8'h9A, 8'h00, 8'hB0, 8'h0A, 8'h69, 8'h04, 8'hD9, 8'h9A, 8'h00, 8'h90, 8'h03,
			8'h20, 8'hBF, 8'hCC, 8'hB9, 8'h91, 8'h00, 8'h18, 8'h69, 8'h08, 8'h38, 8'hFD, 8'hD2, 8'h05, 8'h20, 8'h8E, 8'hF0,
			8'h85, 8'h12, 8'hB9, 8'h9A, 8'h00, 8'h18, 8'h69, 8'h0C, 8'h38, 8'hFD, 8'hDC, 8'h05, 8'h20, 8'h8E, 8'hF0, 8'h85,
			8'h13, 8'hBD, 8'hFA, 8'h05, 8'hC9, 8'h03, 8'hF0, 8'h0A, 8'hA5, 8'h12, 8'h48, 8'hA5, 8'h13, 8'h85, 8'h12, 8'h68,
			8'h85, 8'h13, 8'hA5, 8'h12, 8'hC9, 8'h14, 8'hB0, 8'h10, 8'hA5, 8'h13, 8'hC9, 8'h0B, 8'hB0, 8'h0A, 8'hA9, 8'h01,
			8'h9D, 8'h04, 8'h06, 8'hA9, 8'h32, 8'h9D, 8'h0E, 8'h06, 8'h88, 8'h30, 8'h03, 8'h4C, 8'h3A, 8'hCC, 8'h60, 8'h8A,
			8'h48, 8'h98, 8'hAA, 8'hE6, 8'hCB, 8'h20, 8'h83, 8'hE9, 8'h68, 8'hAA, 8'h60, 8'hBD, 8'hF0, 8'h05, 8'h85, 8'h57,
			8'hBD, 8'hE6, 8'h05, 8'h85, 8'h58, 8'hA9, 8'h03, 8'h85, 8'h59, 8'hBC, 8'hFA, 8'h05, 8'hB9, 8'h26, 8'hCD, 8'h85,
			8'h5A, 8'hB9, 8'h2A, 8'hCD, 8'h85, 8'h5B, 8'hB9, 8'h2E, 8'hCD, 8'h85, 8'h5C, 8'h20, 8'h0F, 8'hCD, 8'hB9, 8'h32,
			8'hCD, 8'h85, 8'h5A, 8'hB9, 8'h36, 8'hCD, 8'h85, 8'h5B, 8'hB9, 8'h3A, 8'hCD, 8'h85, 8'h5C, 8'h20, 8'h0F, 8'hCD,
			8'hB9, 8'h3E, 8'hCD, 8'h85, 8'h5A, 8'hB9, 8'h42, 8'hCD, 8'h85, 8'h5B, 8'hB9, 8'h46, 8'hCD, 8'h85, 8'h5C, 8'h98,
			8'h48, 8'hA9, 8'h57, 8'hA0, 8'h00, 8'h20, 8'h31, 8'hC1, 8'h68, 8'hA8, 8'hA5, 8'h58, 8'h18, 8'h69, 8'h20, 8'h85,
			8'h58, 8'h90, 8'h02, 8'hE6, 8'h57, 8'h60, 8'hA1, 8'h24, 8'h24, 8'h24, 8'hA2, 8'h9E, 8'hAB, 8'h24, 8'h24, 8'h24,
			8'hAC, 8'h24, 8'hA3, 8'h24, 8'hAD, 8'hA8, 8'hA4, 8'h9F, 8'hAE, 8'hA9, 8'hA5, 8'h24, 8'hAF, 8'hAA, 8'h24, 8'h24,
			8'hB0, 8'h24, 8'hA6, 8'hA0, 8'hB1, 8'h24, 8'hA7, 8'h24, 8'h24, 8'h24, 8'hA2, 8'h09, 8'hA9, 8'hFF, 8'h9D, 8'h5D,
			8'h05, 8'hA9, 8'hF0, 8'h9D, 8'h7B, 8'h05, 8'hCA, 8'h10, 8'hF3, 8'h60, 8'hCE, 8'hCC, 8'h05, 8'hF0, 8'h01, 8'h60,
			8'hA5, 8'h1B, 8'h29, 8'h3F, 8'h69, 8'h28, 8'h8D, 8'hCC, 8'h05, 8'hA2, 8'h09, 8'hBD, 8'h5D, 8'h05, 8'h30, 8'h04,
			8'hCA, 8'h10, 8'hF8, 8'h60, 8'hA9, 8'h00, 8'h9D, 8'h5D, 8'h05, 8'h9D, 8'h99, 8'h05, 8'h9D, 8'h8F, 8'h05, 8'hA9,
			8'h80, 8'h9D, 8'h71, 8'h05, 8'h9D, 8'h85, 8'h05, 8'hA9, 8'hD0, 8'h9D, 8'h7B, 8'h05, 8'h20, 8'hB3, 8'hF1, 8'h29,
			8'h03, 8'hA8, 8'hB9, 8'hAE, 8'hCE, 8'h9D, 8'h67, 8'h05, 8'hA0, 8'h00, 8'hA5, 8'h1B, 8'h9D, 8'hB7, 8'h05, 8'h10,
			8'h01, 8'h88, 8'h98, 8'h9D, 8'hC1, 8'h05, 8'hCE, 8'hCB, 8'h05, 8'h60, 8'hA2, 8'h09, 8'hBD, 8'h5D, 8'h05, 8'h30,
			8'h71, 8'hF0, 8'h49, 8'hBD, 8'h99, 8'h05, 8'h85, 8'h12, 8'hBD, 8'h8F, 8'h05, 8'h85, 8'h13, 8'h20, 8'hA6, 8'hF1,
			8'hBD, 8'hB7, 8'h05, 8'h18, 8'h65, 8'h12, 8'h9D, 8'hB7, 8'h05, 8'h85, 8'h12, 8'hBD, 8'hC1, 8'h05, 8'h65, 8'h13,
			8'h9D, 8'hC1, 8'h05, 8'h85, 8'h13, 8'h20, 8'hA6, 8'hF1, 8'hBD, 8'h99, 8'h05, 8'h38, 8'hE5, 8'h12, 8'h9D, 8'h99,
			8'h05, 8'hBD, 8'h8F, 8'h05, 8'hE5, 8'h13, 8'h9D, 8'h8F, 8'h05, 8'hBD, 8'h71, 8'h05, 8'h18, 8'h7D, 8'h99, 8'h05,
			8'h9D, 8'h71, 8'h05, 8'hBD, 8'h67, 8'h05, 8'h7D, 8'h8F, 8'h05, 8'h9D, 8'h67, 8'h05, 8'hBD, 8'h85, 8'h05, 8'h38,
			8'hED, 8'h5A, 8'h05, 8'h9D, 8'h85, 8'h05, 8'hB0, 8'h03, 8'hDE, 8'h7B, 8'h05, 8'hBD, 8'h7B, 8'h05, 8'hC9, 8'hF0,
			8'hF0, 8'h0B, 8'hC9, 8'hA8, 8'hB0, 8'h0C, 8'hA9, 8'h01, 8'h9D, 8'h5D, 8'h05, 8'hD0, 8'h05, 8'hA9, 8'hFF, 8'h9D,
			8'h5D, 8'h05, 8'h20, 8'h2F, 8'hCE, 8'h20, 8'hCE, 8'hCE, 8'hCA, 8'h30, 8'h03, 8'h4C, 8'hAC, 8'hCD, 8'h60, 8'hBC,
			8'h5D, 8'h05, 8'hC8, 8'hB9, 8'hB2, 8'hCE, 8'h85, 8'h13, 8'h8A, 8'h85, 8'h12, 8'h0A, 8'h65, 8'h12, 8'h0A, 8'h0A,
			8'hA8, 8'hBD, 8'h7B, 8'h05, 8'h99, 8'h50, 8'h02, 8'h99, 8'h54, 8'h02, 8'h18, 8'h69, 8'h08, 8'h99, 8'h58, 8'h02,
			8'hBD, 8'h67, 8'h05, 8'h99, 8'h53, 8'h02, 8'h18, 8'h69, 8'h04, 8'h99, 8'h5B, 8'h02, 8'h18, 8'h69, 8'h04, 8'h99,
			8'h57, 8'h02, 8'hA5, 8'h13, 8'h99, 8'h52, 8'h02, 8'h99, 8'h56, 8'h02, 8'h99, 8'h5A, 8'h02, 8'hBD, 8'h5D, 8'h05,
			8'h30, 8'h27, 8'hA9, 8'hA8, 8'h99, 8'h51, 8'h02, 8'hA9, 8'hA9, 8'h99, 8'h55, 8'h02, 8'hA5, 8'h19, 8'h4A, 8'h4A,
			8'h4A, 8'h4A, 8'h29, 8'h07, 8'h86, 8'h13, 8'hAA, 8'hBD, 8'hB5, 8'hCE, 8'h99, 8'h59, 8'h02, 8'hB9, 8'h5A, 8'h02,
			8'h5D, 8'hBD, 8'hCE, 8'h99, 8'h5A, 8'h02, 8'hA6, 8'h13, 8'h60, 8'hA9, 8'hF0, 8'h9D, 8'h7B, 8'h05, 8'hA9, 8'hAC,
			8'h99, 8'h51, 8'h02, 8'hA9, 8'hAD, 8'h99, 8'h55, 8'h02, 8'hA9, 8'hFC, 8'h99, 8'h59, 8'h02, 8'h60, 8'h20, 8'h50,
			8'hA0, 8'hD0, 8'h02, 8'h22, 8'h02, 8'hAA, 8'hAB, 8'hAB, 8'hAA, 8'hAA, 8'hAB, 8'hAB, 8'hAA, 8'h00, 8'h00, 8'h40,
			8'h40, 8'h40, 8'h40, 8'h00, 8'h00, 8'hFC, 8'hFC, 8'hDF, 8'hFC, 8'hFC, 8'hE0, 8'hE2, 8'hE1, 8'hFC, 8'hA0, 8'h01,
			8'hB9, 8'h88, 8'h00, 8'h30, 8'h3A, 8'hF0, 8'h38, 8'hBD, 8'h5D, 8'h05, 8'h30, 8'h36, 8'hB9, 8'h9A, 8'h00, 8'hC9,
			8'hC0, 8'hB0, 8'h2C, 8'h38, 8'hFD, 8'h7B, 8'h05, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h18, 8'hB0, 8'h21, 8'hB9, 8'h91,
			8'h00, 8'h38, 8'hFD, 8'h67, 8'h05, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h10, 8'hB0, 8'h13, 8'hA9, 8'hFF, 8'h9D, 8'h5D,
			8'h05, 8'hB9, 8'hCD, 8'h05, 8'h18, 8'h69, 8'h01, 8'h99, 8'hCD, 8'h05, 8'hA9, 8'h02, 8'h85, 8'hF0, 8'h60, 8'h88,
			8'h10, 8'hBE, 8'h60, 8'hA9, 8'h20, 8'h85, 8'hF2, 8'h20, 8'hE2, 8'hD0, 8'h20, 8'h4A, 8'hCD, 8'hA6, 8'h40, 8'hB5,
			8'h41, 8'h30, 8'h03, 8'h20, 8'hB0, 8'hF3, 8'hCA, 8'h10, 8'hF6, 8'hA2, 8'h00, 8'h86, 8'hBD, 8'h86, 8'hBE, 8'hA9,
			8'h14, 8'h8D, 8'hCB, 8'h05, 8'h20, 8'h70, 8'hF4, 8'hE6, 8'h4C, 8'h20, 8'hDD, 8'hD8, 8'h20, 8'h91, 8'hE6, 8'hAD,
			8'hCB, 8'h05, 8'hF0, 8'h03, 8'h20, 8'h5A, 8'hCD, 8'h20, 8'hAA, 8'hCD, 8'hAD, 8'hCB, 8'h05, 8'hD0, 8'hE5, 8'hA2,
			8'h09, 8'hBD, 8'h5D, 8'h05, 8'h10, 8'hDE, 8'hCA, 8'h10, 8'hF8, 8'hA5, 8'h19, 8'hD0, 8'hD7, 8'h20, 8'h46, 8'hD2,
			8'hA2, 8'h02, 8'h86, 8'h46, 8'h20, 8'h5E, 8'hF4, 8'hA9, 8'h2B, 8'hA0, 8'hD1, 8'h20, 8'h31, 8'hC1, 8'hA9, 8'h5A,
			8'hA0, 8'hD1, 8'h20, 8'h31, 8'hC1, 8'hA9, 8'h65, 8'hA0, 8'hD1, 8'h20, 8'h31, 8'hC1, 8'hA6, 8'h40, 8'hA9, 8'h20,
			8'h95, 8'h91, 8'hBD, 8'h9E, 8'hD1, 8'h95, 8'h9A, 8'hA9, 8'h03, 8'h95, 8'h7F, 8'hA9, 8'h01, 8'h9D, 8'h48, 8'h04,
			8'h20, 8'hB0, 8'hF3, 8'h20, 8'hA4, 8'hE3, 8'hCA, 8'h10, 8'hE5, 8'hA9, 8'h44, 8'h8D, 8'h67, 8'h05, 8'h8D, 8'h68,
			8'h05, 8'hA9, 8'h54, 8'h8D, 8'h7B, 8'h05, 8'hA9, 8'h74, 8'h8D, 8'h7C, 8'h05, 8'hA9, 8'h01, 8'h8D, 8'h5D, 8'h05,
			8'h8D, 8'h5E, 8'h05, 8'hA6, 8'h40, 8'h20, 8'h2F, 8'hCE, 8'hCA, 8'h10, 8'hFA, 8'h20, 8'h5C, 8'hF4, 8'hA9, 8'h2B,
			8'h85, 8'h57, 8'hA9, 8'h24, 8'h85, 8'h58, 8'h85, 8'h59, 8'hA9, 8'h0C, 8'h85, 8'h54, 8'hA9, 8'h0B, 8'h85, 8'h55,
			8'hA9, 8'h05, 8'h85, 8'h56, 8'hAD, 8'hCD, 8'h05, 8'h20, 8'hC9, 8'hD1, 8'hA5, 8'h40, 8'hF0, 8'h0A, 8'hA9, 8'h0F,
			8'h85, 8'h55, 8'hAD, 8'hCE, 8'h05, 8'h20, 8'hC9, 8'hD1, 8'h20, 8'h5C, 8'hF4, 8'hAD, 8'h59, 8'h05, 8'h85, 8'h57,
			8'hA9, 8'h00, 8'h85, 8'h58, 8'h85, 8'h59, 8'hA9, 8'h08, 8'h85, 8'h54, 8'hA9, 8'h0B, 8'h85, 8'h55, 8'hA9, 8'h03,
			8'h85, 8'h56, 8'hAD, 8'h59, 8'h05, 8'h20, 8'h19, 8'hC1, 8'hA5, 8'h40, 8'hF0, 8'h07, 8'hA9, 8'h0F, 8'h85, 8'h55,
			8'h20, 8'h19, 8'hC1, 8'hA9, 8'hFF, 8'h8D, 8'h5D, 8'h05, 8'h8D, 8'h5E, 8'h05, 8'hA6, 8'h40, 8'h20, 8'h2F, 8'hCE,
			8'hCA, 8'h10, 8'hFA, 8'hA9, 8'h02, 8'h85, 8'hF0, 8'hA2, 8'h02, 8'h20, 8'h5E, 8'hF4, 8'hA6, 8'h40, 8'h20, 8'h2F,
			8'hCE, 8'hCA, 8'h10, 8'hFA, 8'h20, 8'hA0, 8'hD1, 8'h20, 8'h5C, 8'hF4, 8'hA9, 8'h01, 8'h85, 8'hF0, 8'h20, 8'h21,
			8'hD1, 8'hD0, 8'h25, 8'hA9, 8'h70, 8'hA0, 8'hD1, 8'h20, 8'h31, 8'hC1, 8'h20, 8'h65, 8'hF4, 8'hA2, 8'h1A, 8'hBD,
			8'h84, 8'hD1, 8'h95, 8'h57, 8'hCA, 8'h10, 8'hF8, 8'hAD, 8'h5B, 8'h05, 8'h85, 8'h68, 8'hAD, 8'h5C, 8'h05, 8'h85,
			8'h69, 8'h20, 8'h2D, 8'hC1, 8'hA9, 8'h10, 8'h85, 8'hF2, 8'hA2, 8'h78, 8'h20, 8'h5E, 8'hF4, 8'h20, 8'hA0, 8'hD1,
			8'hA9, 8'h00, 8'h85, 8'h3E, 8'hA2, 8'h04, 8'h20, 8'h13, 8'hD2, 8'h20, 8'h2D, 8'hC1, 8'hA5, 8'h40, 8'hF0, 8'h0E,
			8'hE6, 8'h3E, 8'hA2, 8'h12, 8'h20, 8'h13, 8'hD2, 8'hA9, 8'h65, 8'hA0, 8'h00, 8'h20, 8'h31, 8'hC1, 8'hA9, 8'h01,
			8'h85, 8'hF1, 8'hA2, 8'h02, 8'h20, 8'h5E, 8'hF4, 8'hA5, 8'h5D, 8'hC9, 8'h24, 8'hD0, 8'hD3, 8'hA5, 8'h40, 8'hF0,
			8'h07, 8'hAD, 8'h6B, 8'h00, 8'hC9, 8'h24, 8'hD0, 8'hC8, 8'hA2, 8'h0A, 8'h20, 8'h5E, 8'hF4, 8'h20, 8'h21, 8'hD1,
			8'hD0, 8'h1C, 8'hAD, 8'h5B, 8'h05, 8'h85, 8'h47, 8'hAD, 8'h5C, 8'h05, 8'h85, 8'h48, 8'hA5, 8'h40, 8'h85, 8'h3E,
			8'h20, 8'hDC, 8'hD6, 8'hC6, 8'h3E, 8'h10, 8'hF9, 8'hA9, 8'h01, 8'h85, 8'hF1, 8'h20, 8'h5C, 8'hF4, 8'hA9, 8'h00,
			8'h85, 8'h47, 8'h85, 8'h48, 8'hA2, 8'h01, 8'hB5, 8'h41, 8'h10, 8'h02, 8'h95, 8'h88, 8'hCA, 8'h10, 8'hF7, 8'h4C,
			8'h53, 8'hF3, 8'hAE, 8'h58, 8'h05, 8'hBD, 8'h0D, 8'hD1, 8'h8D, 8'h59, 8'h05, 8'hBD, 8'h12, 8'hD1, 8'h8D, 8'h5A,
			8'h05, 8'hBD, 8'h17, 8'hD1, 8'h8D, 8'h5B, 8'h05, 8'hBD, 8'h1C, 8'hD1, 8'h8D, 8'h5C, 8'h05, 8'hE0, 8'h04, 8'hB0,
			8'h03, 8'hEE, 8'h58, 8'h05, 8'hA9, 8'h00, 8'h8D, 8'hCD, 8'h05, 8'h8D, 8'hCE, 8'h05, 8'h60, 8'h03, 8'h05, 8'h07,
			8'h07, 8'h07, 8'h80, 8'h90, 8'h98, 8'hA0, 8'hA8, 8'h01, 8'h01, 8'h02, 8'h02, 8'h03, 8'h00, 8'h05, 8'h00, 8'h05,
			8'h00, 8'hAD, 8'hCD, 8'h05, 8'h18, 8'h6D, 8'hCE, 8'h05, 8'hC9, 8'h14, 8'h60, 8'h3F, 8'h00, 8'h10, 8'h0F, 8'h30,
			8'h30, 8'h30, 8'h0F, 8'h30, 8'h27, 8'h15, 8'h0F, 8'h30, 8'h02, 8'h21, 8'h0F, 8'h16, 8'h16, 8'h16, 8'h21, 8'h73,
			8'h0B, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h19, 8'h1D, 8'h1C, 8'h26, 8'h21, 8'hF3, 8'h0B, 8'h29,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h19, 8'h1D, 8'h1C, 8'h26, 8'h23, 8'hE8, 8'h08, 8'hFF, 8'hFF, 8'hFF,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h23, 8'hC0, 8'h08, 8'h40, 8'h50, 8'h50, 8'h50, 8'h50, 8'h90, 8'hA0, 8'hA0,
			8'h22, 8'h88, 8'h11, 8'h19, 8'h24, 8'h0E, 8'h24, 8'h1B, 8'h24, 8'h0F, 8'h24, 8'h0E, 8'h24, 8'h0C, 8'h24, 8'h1D,
			8'h24, 8'h2C, 8'h2C, 8'h2C, 8'h22, 8'hC6, 8'h17, 8'h1C, 8'h1E, 8'h19, 8'h0E, 8'h1B, 8'h24, 8'h0B, 8'h18, 8'h17,
			8'h1E, 8'h1C, 8'h24, 8'h24, 8'h24, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h19, 8'h1D, 8'h1C, 8'h2C, 8'h50, 8'h70,
			8'hA2, 8'h1C, 8'hBD, 8'h3E, 8'hD1, 8'h95, 8'h57, 8'hCA, 8'h10, 8'hF8, 8'hA2, 8'h04, 8'hAC, 8'hCD, 8'h05, 8'h20,
			8'hDC, 8'hD1, 8'hA2, 8'h12, 8'hAC, 8'hCE, 8'h05, 8'h20, 8'hDC, 8'hD1, 8'h20, 8'h2D, 8'hC1, 8'hA5, 8'h40, 8'hD0,
			8'h01, 8'h60, 8'hA9, 8'h65, 8'hA0, 8'h00, 8'h4C, 8'h31, 8'hC1, 8'hA0, 8'h00, 8'hC9, 8'h0A, 8'h90, 8'h06, 8'hC8,
			8'hE9, 8'h0A, 8'h4C, 8'hCB, 8'hD1, 8'h84, 8'h5A, 8'h85, 8'h5B, 8'h4C, 8'h19, 8'hC1, 8'h88, 8'h30, 8'h1F, 8'hAD,
			8'h59, 8'h05, 8'h18, 8'h75, 8'h59, 8'hC9, 8'h0A, 8'h90, 8'h04, 8'hE9, 8'h0A, 8'hF6, 8'h58, 8'h95, 8'h59, 8'hB5,
			8'h58, 8'hC9, 8'h0A, 8'h90, 8'h06, 8'hE9, 8'h0A, 8'hF6, 8'h57, 8'h95, 8'h58, 8'h4C, 8'hDC, 8'hD1, 8'hA0, 8'h00,
			8'hB5, 8'h57, 8'hF0, 8'h04, 8'hC9, 8'h24, 8'hD0, 8'h0A, 8'hA9, 8'h24, 8'h95, 8'h57, 8'hE8, 8'hC8, 8'hC0, 8'h04,
			8'hD0, 8'hEE, 8'h60, 8'hB5, 8'h59, 8'hC9, 8'h24, 8'hF0, 8'h2A, 8'hA8, 8'hD0, 8'h1C, 8'hB5, 8'h58, 8'hC9, 8'h24,
			8'hF0, 8'h21, 8'hB5, 8'h58, 8'hD0, 8'h0C, 8'hB5, 8'h57, 8'hC9, 8'h24, 8'hF0, 8'h17, 8'hA9, 8'h0A, 8'h95, 8'h58,
			8'hD6, 8'h57, 8'hA9, 8'h0A, 8'h95, 8'h59, 8'hD6, 8'h58, 8'hD6, 8'h59, 8'h8A, 8'h48, 8'hA9, 8'h0A, 8'h20, 8'hDE,
			8'hD6, 8'h68, 8'hAA, 8'h4C, 8'hFE, 8'hD1, 8'h20, 8'h0A, 8'hC1, 8'h20, 8'hFA, 8'hC0, 8'hA9, 8'h20, 8'h8D, 8'h06,
			8'h20, 8'hA9, 8'h00, 8'h8D, 8'h06, 8'h20, 8'h20, 8'h75, 8'hD2, 8'h20, 8'h75, 8'hD2, 8'h20, 8'h04, 8'hC1, 8'h20,
			8'h15, 8'hC1, 8'hA2, 8'h3F, 8'hA0, 8'h00, 8'h84, 8'h4C, 8'hA9, 8'hF0, 8'h99, 8'h00, 8'h02, 8'hC8, 8'hC8, 8'hC8,
			8'hC8, 8'hCA, 8'h10, 8'hF4, 8'h60, 8'hA2, 8'hF0, 8'hA9, 8'h24, 8'h8D, 8'h07, 8'h20, 8'h8D, 8'h07, 8'h20, 8'h8D,
			8'h07, 8'h20, 8'h8D, 8'h07, 8'h20, 8'hCA, 8'hD0, 8'hF1, 8'hA2, 8'h40, 8'hA9, 8'h00, 8'h8D, 8'h07, 8'h20, 8'hCA,
			8'hD0, 8'hFA, 8'h60, 8'h20, 8'h0A, 8'hC1, 8'h20, 8'hFA, 8'hC0, 8'hA5, 8'h16, 8'hF0, 8'h03, 8'h4C, 8'h72, 8'hD5,
			8'hA4, 8'h3B, 8'hB9, 8'h2A, 8'hDB, 8'h85, 8'h1D, 8'hB9, 8'h3A, 8'hDB, 8'h85, 8'h1E, 8'h20, 8'h97, 8'hD4, 8'hA2,
			8'h00, 8'h20, 8'hE5, 8'hD4, 8'hC9, 8'hFF, 8'hF0, 8'h6A, 8'h85, 8'h54, 8'h20, 8'hE5, 8'hD4, 8'h85, 8'h55, 8'hA0,
			8'h03, 8'h20, 8'hFB, 8'hD4, 8'hA9, 8'h04, 8'h85, 8'h12, 8'hB9, 8'h93, 8'hD4, 8'h8D, 8'h07, 8'h20, 8'h18, 8'h69,
			8'h04, 8'hC6, 8'h12, 8'hD0, 8'hF6, 8'hE6, 8'h55, 8'h88, 8'h10, 8'hE7, 8'hA5, 8'h55, 8'h38, 8'hE9, 8'h04, 8'h85,
			8'h55, 8'h20, 8'h1C, 8'hD5, 8'h95, 8'hA6, 8'hE6, 8'h54, 8'hE6, 8'h54, 8'h20, 8'h1C, 8'hD5, 8'h95, 8'hA9, 8'hE6,
			8'h55, 8'hE6, 8'h55, 8'h20, 8'h1C, 8'hD5, 8'h95, 8'hAF, 8'hC6, 8'h54, 8'hC6, 8'h54, 8'h20, 8'h1C, 8'hD5, 8'h95,
			8'hAC, 8'h86, 8'hA4, 8'hA9, 8'h03, 8'h20, 8'h56, 8'hC8, 8'h20, 8'h7C, 8'hC1, 8'hA6, 8'hA4, 8'hA5, 8'h54, 8'h0A,
			8'h0A, 8'h0A, 8'h18, 8'h69, 8'h10, 8'h95, 8'hB2, 8'hA5, 8'h55, 8'h0A, 8'h0A, 8'h0A, 8'h95, 8'hB5, 8'hE8, 8'h4C,
			8'hB1, 8'hD2, 8'hCA, 8'h86, 8'hA3, 8'hA2, 8'h00, 8'h20, 8'hE5, 8'hD4, 8'hC9, 8'hFF, 8'hF0, 8'h50, 8'h85, 8'h54,
			8'h20, 8'hE5, 8'hD4, 8'h85, 8'h55, 8'h20, 8'hE5, 8'hD4, 8'h9D, 8'hFA, 8'h05, 8'hA5, 8'h54, 8'h0A, 8'h0A, 8'h0A,
			8'h69, 8'h0C, 8'h9D, 8'hD2, 8'h05, 8'hA5, 8'h55, 8'h0A, 8'h0A, 8'h0A, 8'h69, 8'h0C, 8'h9D, 8'hDC, 8'h05, 8'hA9,
			8'h00, 8'h9D, 8'h04, 8'h06, 8'h20, 8'hFB, 8'hD4, 8'h9D, 8'hE6, 8'h05, 8'hA5, 8'h13, 8'h9D, 8'hF0, 8'h05, 8'h20,
			8'h6C, 8'hD5, 8'h20, 8'h3C, 8'hD5, 8'hE6, 8'h54, 8'hE6, 8'h54, 8'h20, 8'h3C, 8'hD5, 8'hE6, 8'h55, 8'hE6, 8'h55,
			8'h20, 8'h3C, 8'hD5, 8'hC6, 8'h54, 8'hC6, 8'h54, 8'h20, 8'h3C, 8'hD5, 8'hE8, 8'h4C, 8'h27, 8'hD3, 8'hCA, 8'h8E,
			8'hD1, 8'h05, 8'h20, 8'hE5, 8'hD4, 8'h85, 8'h1F, 8'h20, 8'hE5, 8'hD4, 8'h85, 8'h20, 8'hA0, 8'h00, 8'hB1, 8'h1F,
			8'hAA, 8'hCA, 8'h10, 8'h05, 8'hE6, 8'hC8, 8'h4C, 8'hBA, 8'hD3, 8'hC8, 8'hB1, 8'h1F, 8'hC8, 8'h95, 8'h93, 8'hB1,
			8'h1F, 8'hC8, 8'h95, 8'h9C, 8'hB1, 8'h1F, 8'hC8, 8'h9D, 8'h53, 8'h04, 8'hA9, 8'h02, 8'h95, 8'h81, 8'hA9, 8'h01,
			8'h95, 8'h8A, 8'hA5, 8'hC6, 8'h9D, 8'h41, 8'h04, 8'hCA, 8'h10, 8'hE0, 8'h20, 8'hE5, 8'hD4, 8'h85, 8'hCD, 8'h20,
			8'hE5, 8'hD4, 8'h85, 8'h23, 8'h20, 8'hE5, 8'hD4, 8'hA8, 8'h85, 8'h24, 8'hA5, 8'h23, 8'h20, 8'h8C, 8'hD4, 8'h85,
			8'h25, 8'h84, 8'h26, 8'h20, 8'h8C, 8'hD4, 8'h85, 8'h27, 8'h84, 8'h28, 8'h20, 8'h8C, 8'hD4, 8'h85, 8'h29, 8'h84,
			8'h2A, 8'h20, 8'hD9, 8'hD5, 8'h20, 8'hED, 8'hD3, 8'h20, 8'h04, 8'hC1, 8'h4C, 8'h15, 8'hC1, 8'hA2, 8'h22, 8'hBD,
			8'h37, 8'hD4, 8'h95, 8'h57, 8'hCA, 8'h10, 8'hF8, 8'hA5, 8'hC8, 8'hD0, 8'h15, 8'hA5, 8'h3B, 8'h29, 8'h0C, 8'h09,
			8'h03, 8'hA8, 8'hA2, 8'h03, 8'hB9, 8'h5A, 8'hD4, 8'h95, 8'h5A, 8'h88, 8'hCA, 8'h10, 8'hF7, 8'h4C, 8'h2D, 8'hC1,
			8'hAE, 8'h58, 8'h05, 8'hBD, 8'h6A, 8'hD4, 8'h85, 8'h1D, 8'hBD, 8'h6F, 8'hD4, 8'h85, 8'h1E, 8'hA2, 8'h03, 8'hA0,
			8'h07, 8'hB1, 8'h1D, 8'h95, 8'h72, 8'h88, 8'hCA, 8'h10, 8'hF8, 8'hA5, 8'h16, 8'hD0, 8'hE0, 8'hB1, 8'h1D, 8'h99,
			8'h5A, 8'h00, 8'h88, 8'h10, 8'hF8, 8'h30, 8'hD6, 8'h3F, 8'h00, 8'h20, 8'h0F, 8'h2A, 8'h09, 8'h07, 8'h0F, 8'h30,
			8'h27, 8'h15, 8'h0F, 8'h30, 8'h02, 8'h21, 8'h0F, 8'h30, 8'h00, 8'h10, 8'h0F, 8'h16, 8'h12, 8'h37, 8'h0F, 8'h12,
			8'h16, 8'h37, 8'h0F, 8'h17, 8'h11, 8'h35, 8'h0F, 8'h17, 8'h11, 8'h2B, 8'h0F, 8'h2A, 8'h09, 8'h07, 8'h0F, 8'h26,
			8'h06, 8'h07, 8'h0F, 8'h1B, 8'h0C, 8'h07, 8'h0F, 8'h2C, 8'h01, 8'h06, 8'h74, 8'h7C, 8'h84, 8'h84, 8'h84, 8'hD4,
			8'hD4, 8'hD4, 8'hD4, 8'hD4, 8'h0F, 8'h02, 8'h08, 8'h06, 8'h0F, 8'h2B, 8'h30, 8'h12, 8'h0F, 8'h07, 8'h0A, 8'h19,
			8'h0F, 8'h26, 8'h30, 8'h2B, 8'h0F, 8'h07, 8'h0C, 8'h1C, 8'h0F, 8'h15, 8'h30, 8'h26, 8'h38, 8'h65, 8'hCD, 8'h90,
			8'h01, 8'hC8, 8'h60, 8'h7F, 8'h7E, 8'h7D, 8'h7C, 8'h20, 8'hE5, 8'hD4, 8'h85, 8'h1F, 8'h20, 8'hE5, 8'hD4, 8'h85,
			8'h20, 8'hAA, 8'hF0, 8'h40, 8'h20, 8'hF0, 8'hD4, 8'hAA, 8'hF0, 8'hED, 8'h29, 8'h7F, 8'h8D, 8'h06, 8'h20, 8'h20,
			8'hF0, 8'hD4, 8'h8D, 8'h06, 8'h20, 8'h20, 8'hF0, 8'hD4, 8'h85, 8'h12, 8'h8A, 8'h29, 8'h80, 8'h4A, 8'h4A, 8'h4A,
			8'h4A, 8'h4A, 8'h05, 8'h00, 8'h8D, 8'h00, 8'h20, 8'h8A, 8'h29, 8'h40, 8'hD0, 8'h0C, 8'h20, 8'hF0, 8'hD4, 8'h8D,
			8'h07, 8'h20, 8'hC6, 8'h12, 8'hD0, 8'hF6, 8'hF0, 8'hCC, 8'h20, 8'hF0, 8'hD4, 8'h8D, 8'h07, 8'h20, 8'hC6, 8'h12,
			8'hD0, 8'hF9, 8'hF0, 8'hC0, 8'h60, 8'hA0, 8'h00, 8'hB1, 8'h1D, 8'hE6, 8'h1D, 8'hD0, 8'h02, 8'hE6, 8'h1E, 8'h60,
			8'hA0, 8'h00, 8'hB1, 8'h1F, 8'hE6, 8'h1F, 8'hD0, 8'h02, 8'hE6, 8'h20, 8'h60, 8'hA5, 8'h55, 8'h85, 8'h12, 8'hA9,
			8'h00, 8'h06, 8'h12, 8'h06, 8'h12, 8'h06, 8'h12, 8'h06, 8'h12, 8'h2A, 8'h06, 8'h12, 8'h2A, 8'h09, 8'h20, 8'h8D,
			8'h06, 8'h20, 8'h85, 8'h13, 8'hA5, 8'h12, 8'h05, 8'h54, 8'h8D, 8'h06, 8'h20, 8'h60, 8'hA5, 8'h55, 8'h29, 8'hFC,
			8'h0A, 8'h85, 8'h12, 8'hA5, 8'h54, 8'h4A, 8'h4A, 8'h05, 8'h12, 8'h09, 8'hC0, 8'h48, 8'hA5, 8'h55, 8'h29, 8'h02,
			8'h85, 8'h12, 8'hA5, 8'h54, 8'h29, 8'h02, 8'h4A, 8'h05, 8'h12, 8'hA8, 8'h68, 8'h60, 8'hA9, 8'h23, 8'h8D, 8'h06,
			8'h20, 8'h20, 8'h1C, 8'hD5, 8'h8D, 8'h06, 8'h20, 8'hAD, 8'h07, 8'h20, 8'hAD, 8'h07, 8'h20, 8'h39, 8'h64, 8'hD5,
			8'h19, 8'h68, 8'hD5, 8'h48, 8'hA9, 8'h23, 8'h8D, 8'h06, 8'h20, 8'h20, 8'h1C, 8'hD5, 8'h8D, 8'h06, 8'h20, 8'h68,
			8'h8D, 8'h07, 8'h20, 8'h60, 8'hFC, 8'hF3, 8'hCF, 8'h3F, 8'h01, 8'h04, 8'h10, 8'h40, 8'h20, 8'hCB, 8'hCC, 8'h4C,
			8'h7C, 8'hC1, 8'hA9, 8'hC0, 8'hA0, 8'h23, 8'h20, 8'h93, 8'hD5, 8'hA9, 8'hC0, 8'hA0, 8'h27, 8'h20, 8'h93, 8'hD5,
			8'hA0, 8'h23, 8'hA9, 8'h60, 8'h20, 8'hB8, 8'hD5, 8'hA0, 8'h27, 8'hA9, 8'h60, 8'h20, 8'hB8, 8'hD5, 8'hE6, 8'hC8,
			8'h4C, 8'hE1, 8'hD3, 8'h8C, 8'h06, 8'h20, 8'h8D, 8'h06, 8'h20, 8'hA2, 8'h00, 8'hBD, 8'hAE, 8'hDC, 8'h8D, 8'h07,
			8'h20, 8'hE8, 8'hE0, 8'h08, 8'hD0, 8'hF5, 8'hA9, 8'h00, 8'hA2, 8'h28, 8'h20, 8'hB1, 8'hD5, 8'hA9, 8'hAA, 8'hA2,
			8'h10, 8'h8D, 8'h07, 8'h20, 8'hCA, 8'hD0, 8'hFA, 8'h60, 8'h8C, 8'h06, 8'h20, 8'h8D, 8'h06, 8'h20, 8'hA2, 8'h20,
			8'hA9, 8'h58, 8'h20, 8'hC9, 8'hD5, 8'hA2, 8'h40, 8'hA9, 8'h5C, 8'h85, 8'h12, 8'h8A, 8'h29, 8'h03, 8'h49, 8'h03,
			8'h05, 8'h12, 8'h8D, 8'h07, 8'h20, 8'hCA, 8'hD0, 8'hF3, 8'h60, 8'hA2, 8'h00, 8'h20, 8'h51, 8'hD6, 8'h20, 8'hF1,
			8'hD5, 8'hA5, 8'h51, 8'h09, 8'h04, 8'h85, 8'h51, 8'h20, 8'hF1, 8'hD5, 8'hE8, 8'hE8, 8'hE0, 8'h80, 8'hD0, 8'hEB,
			8'h60, 8'hA5, 8'h51, 8'h8D, 8'h06, 8'h20, 8'hA5, 8'h50, 8'h8D, 8'h06, 8'h20, 8'hAD, 8'h07, 8'h20, 8'hAD, 8'h07,
			8'h20, 8'hC9, 8'h24, 8'hD0, 8'h07, 8'h8A, 8'h29, 8'h03, 8'hA8, 8'h4C, 8'h3B, 8'hD6, 8'h60, 8'hA5, 8'h4C, 8'hF0,
			8'h29, 8'hC6, 8'h4C, 8'hA5, 8'h4F, 8'h18, 8'h69, 8'h02, 8'h29, 8'h3F, 8'h85, 8'h4F, 8'hAA, 8'h20, 8'h51, 8'hD6,
			8'hA5, 8'h51, 8'h8D, 8'h06, 8'h20, 8'hA5, 8'h50, 8'h8D, 8'h06, 8'h20, 8'hAD, 8'h07, 8'h20, 8'hAD, 8'h07, 8'h20,
			8'hA0, 8'h03, 8'hD9, 8'h4C, 8'hD6, 8'hF0, 8'h04, 8'h88, 8'h10, 8'hF8, 8'h60, 8'hA5, 8'h51, 8'h8D, 8'h06, 8'h20,
			8'hA5, 8'h50, 8'h8D, 8'h06, 8'h20, 8'hB9, 8'h4D, 8'hD6, 8'h8D, 8'h07, 8'h20, 8'h60, 8'h24, 8'hED, 8'hEE, 8'hEF,
			8'h24, 8'hBD, 8'h5C, 8'hD6, 8'h85, 8'h50, 8'hBD, 8'h5D, 8'hD6, 8'h85, 8'h51, 8'h60, 8'h63, 8'h21, 8'hA5, 8'h21,
			8'hCB, 8'h20, 8'hB7, 8'h20, 8'h7D, 8'h21, 8'h9B, 8'h22, 8'hF2, 8'h20, 8'h49, 8'h22, 8'h6D, 8'h21, 8'h0B, 8'h22,
			8'h92, 8'h22, 8'h95, 8'h21, 8'h1C, 8'h21, 8'h48, 8'h21, 8'hE0, 8'h20, 8'h0B, 8'h23, 8'hCE, 8'h20, 8'hD0, 8'h21,
			8'h06, 8'h21, 8'h19, 8'h21, 8'h30, 8'h22, 8'h8A, 8'h22, 8'h88, 8'h22, 8'hA4, 8'h20, 8'h42, 8'h22, 8'h68, 8'h21,
			8'h3C, 8'h22, 8'h36, 8'h21, 8'hCA, 8'h21, 8'hBC, 8'h20, 8'h96, 8'h21, 8'h4C, 8'h21, 8'h35, 8'h22, 8'hEF, 8'h20,
			8'h68, 8'h22, 8'hA6, 8'h20, 8'hBB, 8'h21, 8'h7A, 8'h21, 8'hEA, 8'h20, 8'hF1, 8'h21, 8'hC2, 8'h20, 8'h77, 8'h21,
			8'h54, 8'h21, 8'hBA, 8'h20, 8'hC5, 8'h22, 8'hBE, 8'h20, 8'hFA, 8'h20, 8'hAE, 8'h21, 8'h46, 8'h21, 8'h9A, 8'h21,
			8'hD2, 8'h20, 8'h3D, 8'h21, 8'h2B, 8'h22, 8'hB0, 8'h20, 8'hB6, 8'h21, 8'hAC, 8'h20, 8'hB3, 8'h20, 8'hDB, 8'h20,
			8'hF6, 8'h20, 8'h2C, 8'h21, 8'hE7, 8'h20, 8'h62, 8'h21, 8'hE4, 8'h21, 8'h4E, 8'h21, 8'hA9, 8'h00, 8'h85, 8'h43,
			8'hA5, 8'h3A, 8'hF0, 8'h01, 8'h60, 8'hA6, 8'h3E, 8'hE0, 8'h02, 8'hB0, 8'hF9, 8'hB5, 8'h41, 8'h30, 8'hF5, 8'hA0,
			8'h64, 8'h20, 8'h7C, 8'hD7, 8'h18, 8'h65, 8'h48, 8'h85, 8'h45, 8'hA0, 8'h0A, 8'h20, 8'h7C, 8'hD7, 8'h85, 8'h44,
			8'hA6, 8'h3F, 8'hBD, 8'h79, 8'hD7, 8'h85, 8'h21, 8'hA9, 8'h06, 8'h85, 8'h22, 8'hA5, 8'h3E, 8'h0A, 8'h0A, 8'h05,
			8'h3E, 8'hAA, 8'h18, 8'hB5, 8'h03, 8'h65, 8'h43, 8'h20, 8'h8F, 8'hD7, 8'h95, 8'h03, 8'hB5, 8'h04, 8'h65, 8'h44,
			8'h20, 8'h8F, 8'hD7, 8'h95, 8'h04, 8'hB5, 8'h05, 8'h65, 8'h45, 8'h20, 8'h8F, 8'hD7, 8'h95, 8'h05, 8'hB5, 8'h06,
			8'h65, 8'h47, 8'h20, 8'h8F, 8'hD7, 8'h95, 8'h06, 8'hB5, 8'h07, 8'h69, 8'h00, 8'h20, 8'h8F, 8'hD7, 8'h95, 8'h07,
			8'hE8, 8'hE8, 8'hE8, 8'hE8, 8'hA0, 8'h04, 8'hB5, 8'h03, 8'hD1, 8'h21, 8'h90, 8'h19, 8'hD0, 8'h04, 8'hCA, 8'h88,
			8'h10, 8'hF4, 8'hA0, 8'h00, 8'hA5, 8'h3E, 8'h0A, 8'h0A, 8'h05, 8'h3E, 8'hAA, 8'hB5, 8'h03, 8'h91, 8'h21, 8'hE8,
			8'hC8, 8'hC0, 8'h05, 8'hD0, 8'hF6, 8'hA0, 8'h04, 8'hB1, 8'h21, 8'h99, 8'h0D, 8'h00, 8'h88, 8'h10, 8'hF8, 8'hE6,
			8'h46, 8'hA5, 8'h16, 8'hF0, 8'h03, 8'h20, 8'h39, 8'hC5, 8'h60, 8'h29, 8'h2E, 8'h33, 8'h84, 8'h12, 8'hA2, 8'hFF,
			8'hA5, 8'h43, 8'h38, 8'hE5, 8'h12, 8'hE8, 8'hB0, 8'hFA, 8'h18, 8'h65, 8'h12, 8'h85, 8'h43, 8'h8A, 8'h60, 8'hC9,
			8'h0A, 8'hB0, 8'h01, 8'h60, 8'h38, 8'hE9, 8'h0A, 8'h60, 8'hA4, 8'h46, 8'h88, 8'hF0, 8'h03, 8'h10, 8'h66, 8'h60,
			8'hA9, 8'h20, 8'h8D, 8'h06, 8'h20, 8'hA9, 8'h43, 8'h8D, 8'h06, 8'h20, 8'hA9, 8'h8E, 8'h8D, 8'h07, 8'h20, 8'hA2,
			8'h04, 8'hB5, 8'h03, 8'h8D, 8'h07, 8'h20, 8'hCA, 8'h10, 8'hF8, 8'hA9, 8'h00, 8'h8D, 8'h07, 8'h20, 8'hA9, 8'h24,
			8'h8D, 8'h07, 8'h20, 8'h8D, 8'h07, 8'h20, 8'hA2, 8'h8C, 8'h8E, 8'h07, 8'h20, 8'hE8, 8'h8E, 8'h07, 8'h20, 8'hA2,
			8'h04, 8'hB5, 8'h0D, 8'h8D, 8'h07, 8'h20, 8'hCA, 8'h10, 8'hF8, 8'hA9, 8'h00, 8'h8D, 8'h07, 8'h20, 8'hA9, 8'h24,
			8'h8D, 8'h07, 8'h20, 8'h8D, 8'h07, 8'h20, 8'hA5, 8'h16, 8'hD0, 8'h6A, 8'hA5, 8'h40, 8'hF0, 8'h14, 8'hA9, 8'h8F,
			8'h8D, 8'h07, 8'h20, 8'hA2, 8'h04, 8'hB5, 8'h08, 8'h8D, 8'h07, 8'h20, 8'hCA, 8'h10, 8'hF8, 8'hA9, 8'h00, 8'h8D,
			8'h07, 8'h20, 8'hC6, 8'h46, 8'h60, 8'hC6, 8'h46, 8'hA9, 8'h20, 8'h8D, 8'h06, 8'h20, 8'hA9, 8'h62, 8'h8D, 8'h06,
			8'h20, 8'hA5, 8'h41, 8'h20, 8'h26, 8'hD8, 8'hA5, 8'h40, 8'hF0, 8'h20, 8'hA9, 8'h20, 8'h8D, 8'h06, 8'h20, 8'hA9,
			8'h75, 8'h8D, 8'h06, 8'h20, 8'hA5, 8'h42, 8'h30, 8'h13, 8'h85, 8'h50, 8'hA2, 8'h06, 8'hA9, 8'h24, 8'hE4, 8'h50,
			8'hB0, 8'h02, 8'hA9, 8'h2A, 8'h8D, 8'h07, 8'h20, 8'hCA, 8'h10, 8'hF2, 8'h60, 8'hA5, 8'h40, 8'hF0, 8'hE9, 8'hA2,
			8'h08, 8'hBD, 8'h4B, 8'hD8, 8'h8D, 8'h07, 8'h20, 8'hCA, 8'h10, 8'hF7, 8'h60, 8'h1B, 8'h0E, 8'h1F, 8'h18, 8'h24,
			8'h0E, 8'h16, 8'h0A, 8'h10, 8'hA0, 8'h04, 8'hB9, 8'h6C, 8'hD8, 8'h8D, 8'h07, 8'h20, 8'h88, 8'h10, 8'hF7, 8'hA5,
			8'h4A, 8'h8D, 8'h07, 8'h20, 8'hA5, 8'h49, 8'h8D, 8'h07, 8'h20, 8'hC6, 8'h46, 8'h60, 8'hFB, 8'hFA, 8'hF9, 8'hF8,
			8'hF7, 8'h85, 8'h12, 8'h86, 8'h13, 8'h84, 8'h14, 8'hA2, 8'h01, 8'hBD, 8'h1A, 8'h06, 8'h30, 8'h0E, 8'hCA, 8'h10,
			8'hF8, 8'hA2, 8'h01, 8'hAD, 8'h19, 8'h06, 8'hCD, 8'h18, 8'h06, 8'h90, 8'h01, 8'hCA, 8'hA9, 8'h64, 8'h9D, 8'h18,
			8'h06, 8'hA5, 8'h12, 8'h9D, 8'h1A, 8'h06, 8'hA8, 8'h8A, 8'h0A, 8'h0A, 8'h0A, 8'hAA, 8'hB9, 8'hD1, 8'hD8, 8'h9D,
			8'hF1, 8'h02, 8'hB9, 8'hD7, 8'hD8, 8'h9D, 8'hF5, 8'h02, 8'hA4, 8'h13, 8'hB9, 8'h9A, 8'h00, 8'h38, 8'hE9, 8'h08,
			8'h9D, 8'hF0, 8'h02, 8'h9D, 8'hF4, 8'h02, 8'hB9, 8'h91, 8'h00, 8'h9D, 8'hF3, 8'h02, 8'h18, 8'h69, 8'h08, 8'h9D,
			8'hF7, 8'h02, 8'hA5, 8'h3E, 8'h9D, 8'hF2, 8'h02, 8'h9D, 8'hF6, 8'h02, 8'hA4, 8'h14, 8'hA6, 8'h13, 8'hA5, 8'h12,
			8'h60, 8'hF4, 8'hF5, 8'hF6, 8'hF7, 8'hF8, 8'hF9, 8'hFB, 8'hFB, 8'hFA, 8'hFB, 8'hFB, 8'hFB, 8'hA2, 8'h01, 8'hBD,
			8'h1A, 8'h06, 8'h30, 8'h17, 8'hDE, 8'h18, 8'h06, 8'hD0, 8'h12, 8'hA9, 8'hFF, 8'h9D, 8'h1A, 8'h06, 8'h8A, 8'h0A,
			8'h0A, 8'h0A, 8'hA8, 8'hA9, 8'hF0, 8'h99, 8'hF0, 8'h02, 8'h99, 8'hF4, 8'h02, 8'hCA, 8'h10, 8'hE1, 8'h60, 8'hA2,
			8'h01, 8'hA9, 8'h00, 8'h9D, 8'h18, 8'h06, 8'hA9, 8'hFF, 8'h9D, 8'h1A, 8'h06, 8'hCA, 8'h10, 8'hF3, 8'h60, 8'h20,
			8'h46, 8'hD2, 8'h20, 8'h0A, 8'hC1, 8'h20, 8'h65, 8'hF4, 8'h20, 8'hFA, 8'hC0, 8'hA9, 8'h2C, 8'h85, 8'h1D, 8'hA9,
			8'hD9, 8'h85, 8'h1E, 8'h20, 8'h97, 8'hD4, 8'h20, 8'h04, 8'hC1, 8'h4C, 8'h15, 8'hC1, 8'h30, 8'hD9, 8'h00, 8'h00,
			8'h3F, 8'h00, 8'h04, 8'h0F, 8'h30, 8'h27, 8'h2A, 8'h3F, 8'h18, 8'h04, 8'h0F, 8'h16, 8'h30, 8'h21, 8'h20, 8'h7C,
			8'h21, 8'hF0, 8'hF1, 8'h24, 8'h24, 8'h24, 8'h24, 8'hE0, 8'hE1, 8'hE1, 8'hE2, 8'hE0, 8'hE1, 8'hE1, 8'hE2, 8'hE0,
			8'hE2, 8'h24, 8'hE0, 8'hE2, 8'h24, 8'hE0, 8'hE1, 8'hE1, 8'hE2, 8'hE0, 8'hE1, 8'hE1, 8'hE2, 8'hE0, 8'hEC, 8'h24,
			8'hE0, 8'hE2, 8'h20, 8'hA2, 8'h1B, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'hE3, 8'hE5, 8'h24,
			8'hE3, 8'hE5, 8'h24, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'hE3, 8'hE3, 8'hF3, 8'hE3, 8'hE5,
			8'h20, 8'hC2, 8'h1B, 8'hE3, 8'hE4, 8'hE3, 8'hE7, 8'hE3, 8'hE4, 8'hE3, 8'hE5, 8'hE3, 8'hE5, 8'h24, 8'hE3, 8'hE5,
			8'h24, 8'hE3, 8'hE4, 8'hE3, 8'hE5, 8'hE3, 8'hE4, 8'hE3, 8'hE5, 8'hE3, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'h20, 8'hE2,
			8'h1B, 8'hE3, 8'hE3, 8'hE3, 8'hE2, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'hE3, 8'hE5, 8'h24, 8'hE3, 8'hE5, 8'h24, 8'hE3,
			8'hE3, 8'hE3, 8'hE5, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'hE3, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'h21, 8'h02, 8'h1B, 8'hE3,
			8'hE4, 8'hE3, 8'hE5, 8'hE3, 8'hF2, 8'hE3, 8'hE5, 8'hE3, 8'hE3, 8'hE2, 8'hE3, 8'hE3, 8'hE2, 8'hE3, 8'hE3, 8'hE3,
			8'hE5, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'hE3, 8'hF2, 8'hE3, 8'hE3, 8'hE5, 8'h21, 8'h22, 8'h1B, 8'hE6, 8'hE3, 8'hE3,
			8'hE7, 8'hEB, 8'h24, 8'hE6, 8'hE7, 8'hE6, 8'hE3, 8'hE7, 8'hE6, 8'hE3, 8'hE7, 8'hE6, 8'hE3, 8'hE3, 8'hE7, 8'hE6,
			8'hE3, 8'hE3, 8'hE7, 8'hEB, 8'h24, 8'hE6, 8'hE3, 8'hE7, 8'h21, 8'h4C, 8'h12, 8'hE0, 8'hE1, 8'hE1, 8'hE2, 8'hE0,
			8'hE2, 8'hE0, 8'hE1, 8'hE1, 8'hE2, 8'hE8, 8'h24, 8'hE0, 8'hE2, 8'hE0, 8'hE1, 8'hE1, 8'hE2, 8'h21, 8'h6C, 8'h12,
			8'hE3, 8'hE3, 8'hE3, 8'hE7, 8'hE3, 8'hE5, 8'hE3, 8'hF5, 8'hF6, 8'hE7, 8'hE3, 8'hF3, 8'hE3, 8'hE5, 8'hE6, 8'hE3,
			8'hE3, 8'hE7, 8'h21, 8'h8C, 8'h12, 8'hE3, 8'hE3, 8'hEF, 8'h24, 8'hE3, 8'hE5, 8'hE3, 8'h24, 8'h24, 8'h24, 8'hE3,
			8'hE3, 8'hE3, 8'hE5, 8'h24, 8'hE3, 8'hE5, 8'h24, 8'h21, 8'hAC, 8'h12, 8'hE3, 8'hE3, 8'hE1, 8'hEA, 8'hE3, 8'hE5,
			8'hE3, 8'hE9, 8'hE3, 8'hE2, 8'hE3, 8'hE3, 8'hE3, 8'hE5, 8'h24, 8'hE3, 8'hE5, 8'h24, 8'h21, 8'hCC, 8'h12, 8'hE3,
			8'hE3, 8'hEF, 8'h24, 8'hE3, 8'hE5, 8'hE3, 8'hF3, 8'hE3, 8'hE5, 8'hE3, 8'hF2, 8'hE3, 8'hE5, 8'h24, 8'hE3, 8'hE5,
			8'h24, 8'h21, 8'hEC, 8'h12, 8'hE6, 8'hE7, 8'h24, 8'h24, 8'hE6, 8'hE7, 8'hE6, 8'hE7, 8'hE6, 8'hE7, 8'hEB, 8'h24,
			8'hE6, 8'hE7, 8'h24, 8'hE6, 8'hE7, 8'h24, 8'h22, 8'h48, 8'h10, 8'h0A, 8'h24, 8'h24, 8'h01, 8'h25, 8'h19, 8'h15,
			8'h0A, 8'h22, 8'h0E, 8'h1B, 8'h24, 8'h10, 8'h0A, 8'h16, 8'h0E, 8'h22, 8'h88, 8'h10, 8'h0B, 8'h24, 8'h24, 8'h02,
			8'h25, 8'h19, 8'h15, 8'h0A, 8'h22, 8'h0E, 8'h1B, 8'h24, 8'h10, 8'h0A, 8'h16, 8'h0E, 8'h22, 8'hC8, 8'h10, 8'h0C,
			8'h24, 8'h24, 8'h0B, 8'h0A, 8'h15, 8'h15, 8'h18, 8'h18, 8'h17, 8'h24, 8'h24, 8'h1D, 8'h1B, 8'h12, 8'h19, 8'h23,
			8'h49, 8'h0E, 8'hF4, 8'h01, 8'h09, 8'h08, 8'h04, 8'h24, 8'h17, 8'h12, 8'h17, 8'h1D, 8'h0E, 8'h17, 8'h0D, 8'h18,
			8'h00, 8'h20, 8'h04, 8'hC1, 8'h20, 8'h0F, 8'hD9, 8'hA9, 8'h00, 8'h85, 8'h19, 8'h20, 8'h65, 8'hF4, 8'hA5, 8'h19,
			8'hF0, 8'h1F, 8'h20, 8'h08, 8'hDB, 8'h20, 8'h68, 8'hE7, 8'hAA, 8'h29, 8'h10, 8'hD0, 8'h13, 8'h8A, 8'h29, 8'h20,
			8'hF0, 8'h0B, 8'hA9, 8'h00, 8'h85, 8'h19, 8'hA6, 8'h3F, 8'hBD, 8'h05, 8'hDB, 8'h85, 8'h3F, 8'h4C, 8'hCB, 8'hDA,
			8'h60, 8'hE6, 8'h3A, 8'hE6, 8'h40, 8'hA9, 8'h00, 8'h8D, 8'h15, 8'h40, 8'h85, 8'h16, 8'h20, 8'hF2, 8'hF1, 8'hA9,
			8'h00, 8'h85, 8'h3A, 8'hF0, 8'hBC, 8'h01, 8'h02, 8'h00, 8'hA5, 8'h3F, 8'h4A, 8'h85, 8'h16, 8'hA5, 8'h3F, 8'hAA,
			8'h29, 8'h01, 8'h85, 8'h40, 8'hBD, 8'h27, 8'hDB, 8'h8D, 8'h7B, 8'h05, 8'hA9, 8'h2C, 8'h8D, 8'h67, 8'h05, 8'hA2,
			8'h00, 8'h8E, 8'h5D, 8'h05, 8'h4C, 8'h2F, 8'hCE, 8'h8C, 8'h9C, 8'hAC, 8'h4A, 8'h59, 8'hF2, 8'h6C, 8'h77, 8'h88,
			8'hE1, 8'h6C, 8'h99, 8'h03, 8'hCA, 8'h6C, 8'hAD, 8'h17, 8'hE1, 8'h6C, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB,
			8'hDB, 8'hDB, 8'hDB, 8'hDC, 8'hDB, 8'hDB, 8'hDB, 8'hDC, 8'hDB, 8'hDB, 8'h2B, 8'hDC, 8'h39, 8'hDD, 8'h00, 8'h00,
			8'h10, 8'h06, 8'hFF, 8'hFF, 8'h96, 8'hDF, 8'h02, 8'h7A, 8'hDE, 8'h2B, 8'hDC, 8'h39, 8'hDD, 8'h4B, 8'hDD, 8'h00,
			8'h00, 8'h18, 8'h0C, 8'h04, 8'h0E, 8'hFF, 8'hFF, 8'hA0, 8'hDF, 8'h04, 8'h86, 8'hDE, 8'hCA, 8'hDC, 8'h00, 8'h00,
			8'hFF, 8'hFF, 8'hB0, 8'hDF, 8'h00, 8'h9A, 8'hDE, 8'h2B, 8'hDC, 8'h5E, 8'hDD, 8'h00, 8'h00, 8'h08, 8'h06, 8'h18,
			8'h0A, 8'hFF, 8'hFF, 8'hB1, 8'hDF, 8'h06, 8'h9E, 8'hDE, 8'h2B, 8'hDC, 8'h7D, 8'hDD, 8'h00, 8'h00, 8'h04, 8'h06,
			8'h12, 8'h08, 8'hFF, 8'hFF, 8'hC1, 8'hDF, 8'h07, 8'hBA, 8'hDE, 8'h2B, 8'hDC, 8'hA3, 8'hDD, 8'h00, 8'h00, 8'h06,
			8'h06, 8'h14, 8'h10, 8'hFF, 8'h0F, 8'h0D, 8'h01, 8'hFF, 8'hD4, 8'hDF, 8'h09, 8'hDA, 8'hDE, 8'h2B, 8'hDC, 8'hCE,
			8'hDD, 8'h00, 8'h00, 8'h04, 8'h06, 8'h10, 8'h0E, 8'hFF, 8'h08, 8'h0E, 8'h03, 8'h0D, 8'h09, 8'h03, 8'h12, 8'h08,
			8'h03, 8'h17, 8'h0D, 8'h03, 8'hFF, 8'hE7, 8'hDF, 8'h03, 8'h02, 8'hDF, 8'h2B, 8'hDC, 8'h5E, 8'hDD, 8'h00, 8'h00,
			8'h10, 8'h06, 8'h1A, 8'h0C, 8'hFF, 8'h08, 8'h08, 8'h01, 8'h18, 8'h04, 8'h01, 8'hFF, 8'hB1, 8'hDF, 8'h06, 8'h9E,
			8'hDE, 8'h2B, 8'hDC, 8'hDB, 8'hDD, 8'h00, 8'h00, 8'h0E, 8'h06, 8'h0C, 8'h14, 8'hFF, 8'hFF, 8'hF7, 8'hDF, 8'h06,
			8'h12, 8'hDF, 8'h2B, 8'hDC, 8'h01, 8'hDE, 8'h00, 8'h00, 8'h04, 8'h08, 8'h16, 8'h10, 8'hFF, 8'hFF, 8'h07, 8'hE0,
			8'h09, 8'h2E, 8'hDF, 8'h2B, 8'hDC, 8'h32, 8'hDE, 8'h00, 8'h00, 8'h04, 8'h10, 8'h18, 8'h10, 8'hFF, 8'h0E, 8'h06,
			8'h01, 8'hFF, 8'h17, 8'hE0, 8'h07, 8'h56, 8'hDF, 8'h2B, 8'hDC, 8'h5B, 8'hDE, 8'h00, 8'h00, 8'h04, 8'h08, 8'h0E,
			8'h10, 8'hFF, 8'h10, 8'h07, 8'h01, 8'hFF, 8'h2A, 8'hE0, 8'h07, 8'h76, 8'hDF, 8'h23, 8'h40, 8'h88, 8'h39, 8'h38,
			8'h39, 8'h38, 8'h39, 8'h38, 8'h39, 8'h33, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24,
			8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h30, 8'h38, 8'h39, 8'h38, 8'h39, 8'h38, 8'h39, 8'h38, 8'h3C, 8'h3B,
			8'h3C, 8'h3B, 8'h3C, 8'h3B, 8'h3C, 8'h3D, 8'h58, 8'h59, 8'h5A, 8'h5B, 8'h58, 8'h59, 8'h5A, 8'h5B, 8'h58, 8'h59,
			8'h5A, 8'h5B, 8'h58, 8'h59, 8'h5A, 8'h5B, 8'h3A, 8'h3B, 8'h3C, 8'h3B, 8'h3C, 8'h3B, 8'h3C, 8'h3B, 8'h60, 8'h61,
			8'h62, 8'h63, 8'h60, 8'h61, 8'h62, 8'h63, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h5C, 8'h5D,
			8'h5E, 8'h5F, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h60, 8'h61, 8'h62, 8'h63, 8'h60, 8'h61, 8'h62, 8'h63, 8'h5C, 8'h5D,
			8'h5E, 8'h5F, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h5C, 8'h5D,
			8'h5E, 8'h5F, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h5C, 8'h5D, 8'h5E, 8'h5F, 8'h40, 8'h50,
			8'h50, 8'h50, 8'h50, 8'h90, 8'hA0, 8'hA0, 8'h23, 8'hF0, 8'h10, 8'h00, 8'h00, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'h00,
			8'h00, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h00, 8'hA3, 8'h04, 8'h04, 8'h93, 8'h94, 8'h94,
			8'h94, 8'hA3, 8'h05, 8'h04, 8'h95, 8'h96, 8'h96, 8'h96, 8'hA2, 8'hEA, 8'h05, 8'h93, 8'h94, 8'h94, 8'h94, 8'h94,
			8'hA2, 8'hEB, 8'h05, 8'h95, 8'h96, 8'h96, 8'h96, 8'h96, 8'hA3, 8'h34, 8'h03, 8'h93, 8'h94, 8'h94, 8'hA3, 8'h35,
			8'h03, 8'h95, 8'h96, 8'h96, 8'hA3, 8'h1A, 8'h04, 8'h93, 8'h94, 8'h94, 8'h94, 8'hA3, 8'h1B, 8'h04, 8'h95, 8'h96,
			8'h96, 8'h96, 8'h63, 8'h80, 8'h20, 8'h97, 8'h23, 8'hA0, 8'h20, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98,
			8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98,
			8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h98, 8'h99, 8'h23, 8'hC0, 8'h08, 8'h40, 8'h50, 8'h50, 8'h50,
			8'h50, 8'h90, 8'hA0, 8'hA0, 8'h63, 8'hE8, 8'h10, 8'hFF, 8'h00, 8'h22, 8'h49, 8'h0E, 8'h30, 8'h31, 8'h32, 8'h31,
			8'h32, 8'h31, 8'h32, 8'h31, 8'h32, 8'h31, 8'h32, 8'h31, 8'h32, 8'h33, 8'h00, 8'h21, 8'h57, 8'h06, 8'h30, 8'h31,
			8'h32, 8'h31, 8'h32, 8'h33, 8'h21, 8'h65, 8'h06, 8'h30, 8'h31, 8'h32, 8'h31, 8'h32, 8'h33, 8'h00, 8'h21, 8'h90,
			8'h03, 8'h30, 8'h31, 8'h33, 8'h22, 8'h26, 8'h03, 8'h30, 8'h31, 8'h33, 8'h22, 8'h57, 8'h03, 8'h30, 8'h31, 8'h33,
			8'h22, 8'h6C, 8'h03, 8'h30, 8'h31, 8'h33, 8'h22, 8'hF2, 8'h03, 8'h30, 8'h31, 8'h33, 8'h00, 8'h20, 8'hCB, 8'h03,
			8'h30, 8'h31, 8'h33, 8'hA1, 8'h6D, 8'h03, 8'h3E, 8'h3F, 8'h40, 8'hA1, 8'h59, 8'h04, 8'h3E, 8'h3F, 8'h3F, 8'h40,
			8'hA1, 8'hA5, 8'h03, 8'h3E, 8'h3F, 8'h40, 8'h22, 8'hAA, 8'h03, 8'h30, 8'h31, 8'h33, 8'h22, 8'hB3, 8'h03, 8'h30,
			8'h31, 8'h33, 8'h00, 8'h20, 8'hE2, 8'h02, 8'h30, 8'h33, 8'h20, 8'hFB, 8'h02, 8'h30, 8'h33, 8'h21, 8'h57, 8'h02,
			8'h30, 8'h33, 8'h21, 8'h93, 8'h02, 8'h30, 8'h33, 8'h22, 8'h0B, 8'h02, 8'h30, 8'h33, 8'h22, 8'h47, 8'h02, 8'h30,
			8'h33, 8'h22, 8'h83, 8'h02, 8'h30, 8'h33, 8'h22, 8'hCF, 8'h04, 8'h30, 8'h31, 8'h32, 8'h33, 8'h00, 8'h22, 8'hCA,
			8'h03, 8'h30, 8'h31, 8'h33, 8'h22, 8'hD2, 8'h03, 8'h30, 8'h31, 8'h33, 8'h00, 8'h21, 8'h08, 8'h04, 8'h30, 8'h31,
			8'h32, 8'h33, 8'h21, 8'h14, 8'h04, 8'h30, 8'h31, 8'h32, 8'h33, 8'hA1, 8'hA5, 8'h04, 8'h3E, 8'h3F, 8'h3F, 8'h40,
			8'hA1, 8'hBA, 8'h04, 8'h3E, 8'h3F, 8'h3F, 8'h40, 8'h22, 8'h6C, 8'h06, 8'h30, 8'h31, 8'h32, 8'h31, 8'h32, 8'h33,
			8'h00, 8'h22, 8'hEE, 8'h04, 8'h30, 8'h31, 8'h32, 8'h33, 8'h20, 8'hF9, 8'h03, 8'h30, 8'h31, 8'h33, 8'hA1, 8'h1A,
			8'h03, 8'h3F, 8'h3F, 8'h40, 8'h21, 8'h90, 8'h03, 8'h30, 8'h31, 8'h33, 8'hA1, 8'hB1, 8'h03, 8'h3F, 8'h3F, 8'h40,
			8'h22, 8'h28, 8'h03, 8'h30, 8'h31, 8'h33, 8'hA2, 8'h49, 8'h03, 8'h3F, 8'h3F, 8'h40, 8'h20, 8'hEA, 8'h02, 8'h30,
			8'h33, 8'h00, 8'hA2, 8'h6C, 8'h03, 8'h3E, 8'h3F, 8'h40, 8'hA2, 8'h73, 8'h03, 8'h3E, 8'h3F, 8'h40, 8'h20, 8'hE4,
			8'h04, 8'h30, 8'h31, 8'h32, 8'h33, 8'h20, 8'hF8, 8'h04, 8'h30, 8'h31, 8'h32, 8'h33, 8'h21, 8'hA8, 8'h04, 8'h30,
			8'h31, 8'h32, 8'h33, 8'h21, 8'hB5, 8'h04, 8'h30, 8'h31, 8'h32, 8'h33, 8'h00, 8'h22, 8'h64, 8'h02, 8'h30, 8'h33,
			8'h22, 8'h08, 8'h02, 8'h30, 8'h33, 8'h21, 8'hAC, 8'h02, 8'h30, 8'h33, 8'h21, 8'hB4, 8'h02, 8'h30, 8'h33, 8'h22,
			8'h18, 8'h02, 8'h30, 8'h33, 8'h22, 8'h7C, 8'h02, 8'h30, 8'h33, 8'h00, 8'h10, 8'hC8, 8'h48, 8'h38, 8'hFF, 8'hB8,
			8'hCF, 8'hCF, 8'h8F, 8'hE0, 8'hE0, 8'h98, 8'h10, 8'hC4, 8'h48, 8'hB8, 8'h28, 8'h3C, 8'hFF, 8'hB8, 8'hE8, 8'h58,
			8'hCF, 8'hCF, 8'h8F, 8'h4F, 8'h57, 8'hE0, 8'hE0, 8'h98, 8'h58, 8'h60, 8'h10, 8'hFF, 8'hDF, 8'hEC, 8'h10, 8'hC8,
			8'h80, 8'h30, 8'hB8, 8'h60, 8'h90, 8'h38, 8'hFF, 8'h98, 8'h48, 8'hD0, 8'h78, 8'hA8, 8'hCF, 8'hCF, 8'h5F, 8'h87,
			8'h8F, 8'h97, 8'hB7, 8'hE0, 8'hE0, 8'h68, 8'h90, 8'h98, 8'hA0, 8'hC0, 8'h10, 8'hC8, 8'h58, 8'h68, 8'hC8, 8'h28,
			8'h50, 8'h98, 8'h38, 8'hFF, 8'h70, 8'h78, 8'hD0, 8'h30, 8'h68, 8'hB0, 8'hCF, 8'hCF, 8'h2F, 8'h57, 8'h4F, 8'h67,
			8'hA7, 8'hA7, 8'hE0, 8'hE0, 8'h38, 8'h6C, 8'h6C, 8'h7C, 8'hB0, 8'hB0, 8'h10, 8'hC8, 8'h12, 8'hDA, 8'hBA, 8'h9A,
			8'h5A, 8'h3A, 8'h1A, 8'h7A, 8'h38, 8'hFF, 8'h1E, 8'hE6, 8'hC6, 8'hA6, 8'h66, 8'h46, 8'h26, 8'h96, 8'hCF, 8'hCF,
			8'h37, 8'h37, 8'h4F, 8'h5F, 8'h7F, 8'h8F, 8'h9F, 8'hAF, 8'hE0, 8'hE0, 8'h40, 8'h40, 8'h58, 8'h68, 8'h88, 8'h98,
			8'hA8, 8'hB8, 8'h10, 8'hC8, 8'h52, 8'h92, 8'h38, 8'hFF, 8'h66, 8'hA6, 8'hCF, 8'hCF, 8'hAF, 8'hAF, 8'hE0, 8'hE0,
			8'hB8, 8'hB8, 8'h10, 8'hC8, 8'h40, 8'hA0, 8'h28, 8'hD0, 8'h60, 8'h38, 8'hFF, 8'h60, 8'hC0, 8'h30, 8'hD8, 8'h90,
			8'hCF, 8'hCF, 8'h3F, 8'h3F, 8'h67, 8'h67, 8'h97, 8'hE0, 8'hE0, 8'h48, 8'h48, 8'h88, 8'h88, 8'hA0, 8'h10, 8'hC8,
			8'h50, 8'hC8, 8'h88, 8'h40, 8'h70, 8'hD0, 8'h88, 8'h48, 8'h38, 8'hFF, 8'h60, 8'hE0, 8'h98, 8'h58, 8'h90, 8'hD8,
			8'h90, 8'h50, 8'hCF, 8'hCF, 8'h37, 8'h37, 8'h5F, 8'h87, 8'hB7, 8'h3C, 8'h64, 8'h8C, 8'hE0, 8'hE0, 8'h40, 8'h40,
			8'h68, 8'h90, 8'hC0, 8'h60, 8'h80, 8'hA8, 8'h10, 8'hC8, 8'h20, 8'hC0, 8'h40, 8'hA8, 8'h60, 8'h98, 8'h38, 8'hFF,
			8'h40, 8'hE0, 8'h60, 8'hC8, 8'h68, 8'hA0, 8'hCF, 8'hCF, 8'h37, 8'h37, 8'h67, 8'h67, 8'h97, 8'h97, 8'hE0, 8'hE0,
			8'h40, 8'h40, 8'h70, 8'h70, 8'hB0, 8'hB0, 8'h10, 8'hC8, 8'h20, 8'h40, 8'h60, 8'hA0, 8'hC0, 8'hE0, 8'h38, 8'hFF,
			8'h30, 8'h50, 8'h70, 8'hB0, 8'hD0, 8'hF0, 8'hCF, 8'hCF, 8'h97, 8'h7F, 8'h67, 8'h67, 8'h7F, 8'h97, 8'hE0, 8'hE0,
			8'hA0, 8'h88, 8'h70, 8'h70, 8'h88, 8'hA0, 8'h03, 8'h58, 8'h78, 8'h04, 8'h78, 8'h78, 8'h04, 8'h98, 8'h78, 8'h04,
			8'h05, 8'hC8, 8'h38, 8'h05, 8'h38, 8'h40, 8'h05, 8'h58, 8'h78, 8'h04, 8'h78, 8'h78, 8'h04, 8'h98, 8'h78, 8'h04,
			8'h00, 8'h05, 8'h94, 8'hA0, 8'h06, 8'h84, 8'h48, 8'h05, 8'h34, 8'h70, 8'h04, 8'h64, 8'h80, 8'h04, 8'hBC, 8'h78,
			8'h04, 8'h06, 8'h5C, 8'h18, 8'h06, 8'h24, 8'h50, 8'h05, 8'h64, 8'h40, 8'h05, 8'hC4, 8'h38, 8'h05, 8'h54, 8'h90,
			8'h04, 8'h9C, 8'h90, 8'h04, 8'h06, 8'h10, 8'h20, 8'h06, 8'hD8, 8'h20, 8'h06, 8'hB8, 8'h38, 8'h05, 8'h98, 8'h48,
			8'h05, 8'h58, 8'h68, 8'h05, 8'h38, 8'h78, 8'h04, 8'h05, 8'h54, 8'h98, 8'h05, 8'h94, 8'h98, 8'h05, 8'h6C, 8'h39,
			8'h06, 8'h94, 8'h31, 8'h06, 8'hBC, 8'h59, 8'h06, 8'h05, 8'h50, 8'h28, 8'h06, 8'hA8, 8'h28, 8'h06, 8'h24, 8'h50,
			8'h06, 8'hCC, 8'h50, 8'h06, 8'h70, 8'h80, 8'h04, 8'h05, 8'h50, 8'h20, 8'h06, 8'hC8, 8'h20, 8'h06, 8'h84, 8'h48,
			8'h05, 8'h44, 8'h70, 8'h05, 8'h78, 8'hA0, 8'h04, 8'h06, 8'h28, 8'h20, 8'h06, 8'hC8, 8'h20, 8'h06, 8'h48, 8'h50,
			8'h05, 8'hB0, 8'h50, 8'h05, 8'h5C, 8'h80, 8'h04, 8'h94, 8'h80, 8'h04, 8'h06, 8'h20, 8'h80, 8'h04, 8'h40, 8'h68,
			8'h05, 8'h60, 8'h50, 8'h06, 8'hA0, 8'h50, 8'h06, 8'hC0, 8'h68, 8'h05, 8'hE0, 8'h80, 8'h04, 8'h08, 8'h08, 8'hF0,
			8'h08, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h08, 8'h08, 8'h00, 8'h00, 8'h01, 8'h08, 8'h08, 8'h09, 8'h00,
			8'h00, 8'hFF, 8'h08, 8'h08, 8'h07, 8'hFE, 8'h00, 8'h00, 8'h06, 8'h08, 8'h08, 8'h02, 8'h00, 8'h00, 8'h0A, 8'h08,
			8'h08, 8'h02, 8'h00, 8'h01, 8'h0A, 8'h08, 8'h09, 8'h04, 8'h00, 8'h00, 8'h0C, 8'h08, 8'h08, 8'h00, 8'h00, 8'hFE,
			8'h08, 8'h08, 8'h06, 8'hFD, 8'hFD, 8'hFD, 8'h05, 8'h05, 8'h05, 8'h08, 8'h08, 8'h08, 8'h00, 8'h00, 8'h00, 8'h08,
			8'h08, 8'h07, 8'h00, 8'h00, 8'hFF, 8'h08, 8'h08, 8'h09, 8'h00, 8'h00, 8'h01, 8'h0A, 8'h08, 8'h08, 8'h02, 8'h00,
			8'h00, 8'h06, 8'h08, 8'h08, 8'hFE, 8'h00, 8'h00, 8'h06, 8'h08, 8'h07, 8'hFE, 8'h00, 8'hFF, 8'h04, 8'h08, 8'h08,
			8'hFC, 8'h00, 8'h00, 8'h08, 8'h08, 8'h0A, 8'h00, 8'h00, 8'h02, 8'h0B, 8'h0B, 8'h0B, 8'h03, 8'h03, 8'h03, 8'h00,
			8'h00, 8'h01, 8'h02, 8'h03, 8'h04, 8'h05, 8'h00, 8'h00, 8'h01, 8'h02, 8'h03, 8'h06, 8'h07, 8'h00, 8'h00, 8'h01,
			8'h02, 8'h03, 8'h06, 8'h08, 8'h00, 8'h09, 8'h0A, 8'h02, 8'h0B, 8'h0C, 8'h05, 8'h00, 8'h00, 8'h01, 8'h02, 8'h03,
			8'h04, 8'h05, 8'h00, 8'h00, 8'h01, 8'h02, 8'h0D, 8'h0E, 8'h05, 8'h00, 8'h1A, 8'h1B, 8'h1C, 8'h1D, 8'h1E, 8'h1F,
			8'h01, 8'h1A, 8'h1B, 8'h20, 8'h1D, 8'h1E, 8'hFC, 8'h00, 8'h1A, 8'h21, 8'h22, 8'h1D, 8'h23, 8'h24, 8'h00, 8'h00,
			8'h38, 8'h35, 8'h0D, 8'h39, 8'h37, 8'h00, 8'h00, 8'h34, 8'h35, 8'h03, 8'h36, 8'h37, 8'h00, 8'h09, 8'h3A, 8'h35,
			8'h0B, 8'h3B, 8'h37, 8'h00, 8'hCE, 8'hCF, 8'hD0, 8'hD1, 8'hD2, 8'hD3, 8'h00, 8'h25, 8'h26, 8'h27, 8'h28, 8'h29,
			8'h2A, 8'h01, 8'h28, 8'h29, 8'h2C, 8'h25, 8'h26, 8'h2B, 8'h00, 8'h4C, 8'hCC, 8'h02, 8'h4D, 8'hCD, 8'h05, 8'h00,
			8'h4C, 8'h2F, 8'h22, 8'h4D, 8'h30, 8'h24, 8'h07, 8'h4C, 8'h2F, 8'h35, 8'h4D, 8'h30, 8'h37, 8'h02, 8'h4C, 8'h2F,
			8'h27, 8'h4D, 8'h30, 8'h2A, 8'h07, 8'h4C, 8'h2F, 8'h2B, 8'h4D, 8'h30, 8'h2C, 8'h00, 8'h0F, 8'h10, 8'h02, 8'h11,
			8'h12, 8'h05, 8'h00, 8'h0F, 8'h10, 8'h02, 8'h11, 8'h19, 8'h07, 8'h00, 8'h0F, 8'h10, 8'h02, 8'h11, 8'h19, 8'h08,
			8'h00, 8'h13, 8'h14, 8'h02, 8'h15, 8'h16, 8'h05, 8'h00, 8'h0F, 8'h10, 8'h02, 8'h11, 8'h12, 8'h05, 8'h03, 8'h13,
			8'h17, 8'h02, 8'h15, 8'h18, 8'h05, 8'h04, 8'h13, 8'h2D, 8'h1C, 8'h15, 8'h2E, 8'h1F, 8'h05, 8'h13, 8'h2D, 8'h20,
			8'h15, 8'h2E, 8'hFC, 8'h04, 8'h13, 8'h2F, 8'h22, 8'h15, 8'h30, 8'h24, 8'h00, 8'h13, 8'h3C, 8'h35, 8'h15, 8'h3D,
			8'h37, 8'h00, 8'h0F, 8'h40, 8'h35, 8'h11, 8'h41, 8'h37, 8'h03, 8'h13, 8'h3E, 8'h35, 8'h15, 8'h3F, 8'h37, 8'h00,
			8'hD4, 8'hD5, 8'hD0, 8'hD6, 8'hD7, 8'hD3, 8'h00, 8'h25, 8'h31, 8'h27, 8'h32, 8'h33, 8'h2A, 8'h02, 8'h25, 8'h31,
			8'h27, 8'h32, 8'h33, 8'h2A, 8'h00, 8'hFC, 8'h48, 8'h42, 8'hFC, 8'h49, 8'h43, 8'h00, 8'hFC, 8'h48, 8'h44, 8'hFC,
			8'h49, 8'h45, 8'h00, 8'hFC, 8'h4A, 8'h46, 8'hFC, 8'h4B, 8'h47, 8'h00, 8'hFC, 8'hA4, 8'hA5, 8'hFC, 8'hA6, 8'hA7,
			8'h08, 8'hFC, 8'h71, 8'hFC, 8'hFC, 8'h72, 8'h73, 8'h08, 8'hFC, 8'h74, 8'hFC, 8'hFC, 8'h75, 8'h76, 8'h08, 8'hFC,
			8'h71, 8'h77, 8'hFC, 8'h72, 8'h73, 8'h08, 8'hFC, 8'h74, 8'h77, 8'hFC, 8'h75, 8'h76, 8'h08, 8'hFC, 8'h71, 8'h78,
			8'hFC, 8'h72, 8'h73, 8'h08, 8'hFC, 8'h74, 8'h78, 8'hFC, 8'h75, 8'h76, 8'h08, 8'hFC, 8'h71, 8'h79, 8'hFC, 8'h72,
			8'h73, 8'h08, 8'hFC, 8'h74, 8'h79, 8'hFC, 8'h75, 8'h76, 8'h00, 8'h4E, 8'h4F, 8'h50, 8'h51, 8'h52, 8'h53, 8'h00,
			8'h4E, 8'h4F, 8'h50, 8'h51, 8'h5E, 8'h58, 8'h00, 8'h4E, 8'h4F, 8'h50, 8'h51, 8'h5E, 8'h5D, 8'h00, 8'h54, 8'h55,
			8'h50, 8'h56, 8'h57, 8'h53, 8'h00, 8'h4E, 8'h4F, 8'h50, 8'h51, 8'h52, 8'h53, 8'h00, 8'h59, 8'h5A, 8'h50, 8'h5B,
			8'h5C, 8'h53, 8'h00, 8'hFC, 8'h5F, 8'h60, 8'hFC, 8'h61, 8'h62, 8'h06, 8'h63, 8'h64, 8'h60, 8'hFC, 8'h65, 8'h62,
			8'h00, 8'h66, 8'h67, 8'h60, 8'h68, 8'h69, 8'h62, 8'h00, 8'h6A, 8'h67, 8'h60, 8'h6B, 8'h69, 8'h62, 8'h00, 8'hFC,
			8'h6C, 8'h6D, 8'hFC, 8'h6E, 8'h6F, 8'h00, 8'hFC, 8'h6C, 8'h6D, 8'hFC, 8'h6E, 8'h70, 8'hAF, 8'hB6, 8'hBD, 8'hB6,
			8'hC4, 8'hCB, 8'hD2, 8'hCB, 8'hD9, 8'hE0, 8'hE7, 8'hE0, 8'hEE, 8'hF5, 8'hFC, 8'hF5, 8'h0A, 8'h0A, 8'h0A, 8'h0A,
			8'h11, 8'h11, 8'h11, 8'h11, 8'h18, 8'h18, 8'h18, 8'h18, 8'h1F, 8'h1F, 8'h1F, 8'h1F, 8'h26, 8'h26, 8'h26, 8'h26,
			8'h2D, 8'h2D, 8'h2D, 8'h2D, 8'h34, 8'h34, 8'h34, 8'h34, 8'h3B, 8'h42, 8'h49, 8'h42, 8'h50, 8'h57, 8'h5E, 8'h57,
			8'h65, 8'h6C, 8'h73, 8'h6C, 8'h7A, 8'h81, 8'h88, 8'h81, 8'h96, 8'h96, 8'h96, 8'h96, 8'h9D, 8'h9D, 8'h9D, 8'h9D,
			8'hA4, 8'hAB, 8'hB2, 8'hAB, 8'hB9, 8'hA4, 8'hB9, 8'hA4, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0,
			8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1,
			8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1,
			8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1,
			8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1,
			8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'h81, 8'h81, 8'h8F, 8'h81, 8'hF5, 8'hF5, 8'h03, 8'hF5, 8'hE1, 8'hE1, 8'hE1, 8'hE1,
			8'hE0, 8'hE0, 8'hE1, 8'hE0, 8'hF8, 8'hFF, 8'h06, 8'hFF, 8'h0D, 8'h14, 8'h1B, 8'h14, 8'h3E, 8'h3E, 8'h22, 8'h29,
			8'h30, 8'h30, 8'h30, 8'h30, 8'hC0, 8'hC0, 8'hC0, 8'hC0, 8'hC0, 8'hC7, 8'hC0, 8'hC7, 8'hCE, 8'hD5, 8'hCE, 8'hD5,
			8'hDC, 8'hE3, 8'hDC, 8'hE3, 8'hEA, 8'hF1, 8'hEA, 8'hF1, 8'h3E, 8'h45, 8'h3E, 8'h45, 8'h37, 8'h37, 8'h37, 8'h37,
			8'hE1, 8'hE1, 8'hE2, 8'hE1, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2,
			8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE1,
			8'hE1, 8'hE1, 8'hE1, 8'hE1, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'hE2, 8'h44, 8'h2C, 8'h00, 8'h00,
			8'h00, 8'h04, 8'h24, 8'h08, 8'h00, 8'h00, 8'hFC, 8'hFC, 8'hFE, 8'hFC, 8'h00, 8'h7B, 8'hFC, 8'hFC, 8'h7C, 8'hFC,
			8'hFC, 8'h00, 8'h7D, 8'h7E, 8'hFC, 8'h7F, 8'h80, 8'hFC, 8'h00, 8'h81, 8'h82, 8'h83, 8'h84, 8'h85, 8'h86, 8'h00,
			8'h87, 8'h88, 8'hFC, 8'h89, 8'h8A, 8'hFC, 8'h00, 8'h8B, 8'h8C, 8'hFC, 8'h8D, 8'h8E, 8'hFC, 8'h00, 8'h8F, 8'h90,
			8'hFC, 8'hFC, 8'hFC, 8'hFC, 8'h55, 8'h5A, 8'h61, 8'h68, 8'h6F, 8'h76, 8'h7D, 8'hE3, 8'hE3, 8'hE3, 8'hE3, 8'hE3,
			8'hE3, 8'hE3, 8'h20, 8'h38, 8'h50, 8'h68, 8'h80, 8'h98, 8'hB0, 8'hC8, 8'h08, 8'h20, 8'h38, 8'hC8, 8'hB0, 8'h98,
			8'h80, 8'h68, 8'h50, 8'h08, 8'hBD, 8'h92, 8'hE3, 8'h85, 8'h1F, 8'hA5, 8'h19, 8'h4A, 8'h90, 8'h05, 8'hBD, 8'h9B,
			8'hE3, 8'h85, 8'h1F, 8'hA9, 8'h02, 8'h85, 8'h20, 8'hB5, 8'h88, 8'h10, 8'h14, 8'hC9, 8'hFF, 8'hF0, 8'h03, 8'h4C,
			8'hD5, 8'hE4, 8'hA0, 8'h14, 8'hA9, 8'hF0, 8'h91, 8'h1F, 8'h88, 8'h88, 8'h88, 8'h88, 8'h10, 8'hF6, 8'h60, 8'hE0,
			8'h08, 8'hF0, 8'h48, 8'hB5, 8'h7F, 8'h0A, 8'h0A, 8'h7D, 8'h36, 8'h04, 8'hE0, 8'h02, 8'hB0, 8'h2A, 8'hB4, 8'h88,
			8'h79, 8'h4C, 8'hE3, 8'hA8, 8'hB9, 8'h4C, 8'hE2, 8'h85, 8'h1D, 8'hB9, 8'h98, 8'hE2, 8'h85, 8'h1E, 8'hB5, 8'hBD,
			8'hF0, 8'h37, 8'hB4, 8'h88, 8'hB9, 8'h4F, 8'hE3, 8'h7D, 8'h36, 8'h04, 8'hA8, 8'hB9, 8'hE4, 8'hE2, 8'h85, 8'h1D,
			8'hB9, 8'hEC, 8'hE2, 8'h85, 8'h1E, 8'h4C, 8'h29, 8'hE4, 8'hB4, 8'h88, 8'h18, 8'h79, 8'h52, 8'hE3, 8'hA8, 8'hB9,
			8'hF4, 8'hE2, 8'h85, 8'h1D, 8'hB9, 8'h20, 8'hE3, 8'h85, 8'h1E, 8'hD0, 8'h0E, 8'hB4, 8'h7F, 8'h30, 8'hA3, 8'hB9,
			8'h84, 8'hE3, 8'h85, 8'h1D, 8'hB9, 8'h8B, 8'hE3, 8'h85, 8'h1E, 8'hB5, 8'h91, 8'h85, 8'h15, 8'hB5, 8'h9A, 8'h85,
			8'h12, 8'h8A, 8'hF0, 8'h10, 8'hE0, 8'h01, 8'hD0, 8'h04, 8'hA9, 8'h01, 8'hD0, 8'h08, 8'hBD, 8'h51, 8'h04, 8'h18,
			8'h69, 8'h02, 8'h29, 8'h03, 8'hBC, 8'h48, 8'h04, 8'hF0, 8'h02, 8'h09, 8'h40, 8'hB4, 8'h88, 8'hC0, 8'h02, 8'hD0,
			8'h08, 8'hB4, 8'h7F, 8'hC0, 8'h05, 8'hD0, 8'h02, 8'h49, 8'h40, 8'hB4, 8'h9A, 8'hC0, 8'hC9, 8'hB0, 8'h04, 8'hE0,
			8'h09, 8'hD0, 8'h02, 8'h09, 8'h20, 8'h85, 8'h14, 8'hA9, 8'h43, 8'h85, 8'h21, 8'hA9, 8'hE0, 8'h85, 8'h22, 8'hBD,
			8'h48, 8'h04, 8'hF0, 8'h08, 8'hA9, 8'h79, 8'h85, 8'h21, 8'hA9, 8'hE0, 8'h85, 8'h22, 8'hA0, 8'h00, 8'hB1, 8'h1D,
			8'hE6, 8'h1D, 8'hD0, 8'h02, 8'hE6, 8'h1E, 8'h0A, 8'h85, 8'h13, 8'h0A, 8'h65, 8'h13, 8'h65, 8'h21, 8'h85, 8'h21,
			8'h90, 8'h02, 8'hE6, 8'h22, 8'h8A, 8'h48, 8'hA2, 8'h05, 8'hA0, 8'h00, 8'hA5, 8'h12, 8'h18, 8'h7D, 8'h3D, 8'hE0,
			8'h91, 8'h1F, 8'h85, 8'h12, 8'hC8, 8'h84, 8'h13, 8'hA0, 8'h00, 8'hB1, 8'h1D, 8'hE6, 8'h1D, 8'hD0, 8'h02, 8'hE6,
			8'h1E, 8'hA4, 8'h13, 8'h91, 8'h1F, 8'hC8, 8'hA5, 8'h14, 8'h91, 8'h1F, 8'hC8, 8'h84, 8'h13, 8'hA0, 8'h00, 8'hA5,
			8'h15, 8'h18, 8'h71, 8'h21, 8'hE6, 8'h21, 8'hD0, 8'h02, 8'hE6, 8'h22, 8'hA4, 8'h13, 8'h91, 8'h1F, 8'hC8, 8'hCA,
			8'h10, 8'hC8, 8'h68, 8'hAA, 8'h60, 8'h8A, 8'h48, 8'hA4, 8'h1F, 8'hB5, 8'h9A, 8'h99, 8'h00, 8'h02, 8'h99, 8'h04,
			8'h02, 8'h18, 8'h69, 8'h08, 8'h99, 8'h08, 8'h02, 8'h99, 8'h0C, 8'h02, 8'hA9, 8'hF0, 8'h99, 8'h10, 8'h02, 8'h99,
			8'h14, 8'h02, 8'hB5, 8'h91, 8'h99, 8'h03, 8'h02, 8'h99, 8'h0B, 8'h02, 8'h18, 8'h69, 8'h08, 8'h99, 8'h07, 8'h02,
			8'h99, 8'h0F, 8'h02, 8'hB5, 8'h9A, 8'hC9, 8'hD0, 8'hA9, 8'h03, 8'h90, 8'h02, 8'hA9, 8'h23, 8'h99, 8'h02, 8'h02,
			8'hB5, 8'h7F, 8'hD0, 8'h3F, 8'hB9, 8'h02, 8'h02, 8'h99, 8'h06, 8'h02, 8'h99, 8'h0A, 8'h02, 8'h99, 8'h0E, 8'h02,
			8'hA9, 8'hDA, 8'h99, 8'h01, 8'h02, 8'hA9, 8'hDB, 8'h99, 8'h05, 8'h02, 8'hA9, 8'hDC, 8'h99, 8'h09, 8'h02, 8'hA9,
			8'hDD, 8'h99, 8'h0D, 8'h02, 8'hA6, 8'h1F, 8'hA5, 8'h19, 8'h29, 8'h20, 8'hF0, 8'h14, 8'hA5, 8'h19, 8'h29, 8'h40,
			8'hD0, 8'h08, 8'hFE, 8'h00, 8'h02, 8'hFE, 8'h04, 8'h02, 8'hD0, 8'h06, 8'hFE, 8'h03, 8'h02, 8'hFE, 8'h0B, 8'h02,
			8'h68, 8'hAA, 8'h60, 8'hB9, 8'h02, 8'h02, 8'h09, 8'h40, 8'h99, 8'h06, 8'h02, 8'h09, 8'h80, 8'h99, 8'h0E, 8'h02,
			8'h29, 8'hBF, 8'h99, 8'h0A, 8'h02, 8'hA9, 8'hDE, 8'h99, 8'h01, 8'h02, 8'h99, 8'h05, 8'h02, 8'h99, 8'h09, 8'h02,
			8'h99, 8'h0D, 8'h02, 8'hDE, 8'h5A, 8'h04, 8'h10, 8'h0C, 8'hA9, 8'hFF, 8'h95, 8'h88, 8'hA9, 8'hF0, 8'h95, 8'h9A,
			8'hA9, 8'h04, 8'h85, 8'hF1, 8'h68, 8'hAA, 8'h60, 8'hA6, 8'hBB, 8'h30, 8'h39, 8'hBD, 8'hC5, 8'hE5, 8'h85, 8'h1D,
			8'hBD, 8'hCA, 8'hE5, 8'h85, 8'h1E, 8'hA0, 8'h00, 8'hA2, 8'h00, 8'hB1, 8'h1D, 8'h9D, 8'hE0, 8'h02, 8'hC8, 8'hE8,
			8'hC9, 8'hF0, 8'hD0, 8'h03, 8'hE8, 8'hE8, 8'hE8, 8'hE0, 8'h10, 8'hD0, 8'hEE, 8'hA0, 8'h0F, 8'hB9, 8'hE0, 8'h02,
			8'h18, 8'h65, 8'hBC, 8'h99, 8'hE0, 8'h02, 8'h88, 8'h88, 8'h88, 8'h88, 8'h10, 8'hF1, 8'hA5, 8'h19, 8'h29, 8'h03,
			8'hD0, 8'h02, 8'hC6, 8'hBB, 8'h60, 8'hFD, 8'hED, 8'hE0, 8'hD6, 8'hCF, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hD0,
			8'hAE, 8'h03, 8'h04, 8'hF0, 8'hF0, 8'hF0, 8'hC8, 8'hAF, 8'h03, 8'h04, 8'hD0, 8'hB0, 8'h03, 8'h04, 8'hF0, 8'hF0,
			8'hC8, 8'hB1, 8'h03, 8'hFC, 8'hC8, 8'hB2, 8'h03, 8'h04, 8'hD0, 8'hB3, 8'h03, 8'h04, 8'hF0, 8'hC8, 8'hB4, 8'h03,
			8'h00, 8'hC8, 8'hB4, 8'h43, 8'h08, 8'hD0, 8'hB5, 8'h03, 8'h00, 8'hD0, 8'hB5, 8'h43, 8'h08, 8'hF0, 8'hF0, 8'hF0,
			8'hF0, 8'h04, 8'h04, 8'h05, 8'h06, 8'h03, 8'h03, 8'h03, 8'h06, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h28, 8'h32, 8'h46,
			8'h78, 8'h00, 8'h00, 8'h00, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0A, 8'h1E, 8'h32, 8'h70, 8'h00, 8'h00, 8'h00,
			8'h70, 8'h00, 8'h00, 8'h00, 8'h00, 8'h14, 8'h3C, 8'h64, 8'hA0, 8'h00, 8'h00, 8'h00, 8'hA0, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h70, 8'hB0, 8'hE0, 8'h40, 8'h80, 8'h80, 8'h80, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h90, 8'h50, 8'h20, 8'hC0, 8'h80, 8'h80, 8'h80,
			8'hC0, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h50, 8'h90, 8'hC0, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h02, 8'h02, 8'h02, 8'h02, 8'hB0, 8'h70, 8'h40, 8'hC0, 8'hC0, 8'hC0, 8'hC0,
			8'hC0, 8'hC0, 8'hC0, 8'hC0, 8'hC0, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'h01, 8'hFE,
			8'hFE, 8'h20, 8'h25, 8'hEE, 8'hA2, 8'h07, 8'hB5, 8'h88, 8'h10, 8'h0A, 8'hC9, 8'hFF, 8'hF0, 8'h44, 8'h20, 8'hBA,
			8'hEC, 8'h4C, 8'hE2, 8'hE6, 8'hE0, 8'h02, 8'h90, 8'h10, 8'hC9, 8'h01, 8'hD0, 8'h0C, 8'hB5, 8'h7F, 8'hC9, 8'h02,
			8'hB0, 8'h06, 8'hA5, 8'hF1, 8'h09, 8'h20, 8'h85, 8'hF1, 8'hDE, 8'h3F, 8'h04, 8'hD0, 8'h1C, 8'hA9, 8'h03, 8'h9D,
			8'h3F, 8'h04, 8'hE0, 8'h02, 8'hB0, 8'h08, 8'hD6, 8'hBF, 8'hD0, 8'h04, 8'hA9, 8'h00, 8'h95, 8'hBD, 8'h20, 8'h18,
			8'hEA, 8'h86, 8'h3E, 8'h20, 8'hC4, 8'hEB, 8'h20, 8'h96, 8'hE7, 8'h20, 8'h58, 8'hEA, 8'h20, 8'h28, 8'hED, 8'h20,
			8'h83, 8'hE9, 8'h20, 8'hA4, 8'hE3, 8'hCA, 8'h10, 8'hAE, 8'h60, 8'hE0, 8'h02, 8'hB0, 8'h18, 8'hA5, 8'h19, 8'h29,
			8'h0F, 8'hD0, 8'h05, 8'h20, 8'hB3, 8'hF1, 8'h95, 8'h31, 8'hA5, 8'h3A, 8'hD0, 8'h09, 8'h20, 8'h6A, 8'hE7, 8'hBD,
			8'h1C, 8'h06, 8'h95, 8'h31, 8'h60, 8'hB5, 8'h9A, 8'hC9, 8'hA0, 8'h90, 8'h07, 8'hB5, 8'h31, 8'h09, 8'h40, 8'h95,
			8'h31, 8'h60, 8'hDE, 8'h5A, 8'h04, 8'hD0, 8'hED, 8'h20, 8'hB3, 8'hF1, 8'hBC, 8'h51, 8'h04, 8'h39, 8'h62, 8'hE7,
			8'h79, 8'h65, 8'hE7, 8'h9D, 8'h5A, 8'h04, 8'h86, 8'h12, 8'hA5, 8'h19, 8'h2A, 8'h2A, 8'h45, 8'h12, 8'h29, 8'h01,
			8'hA8, 8'hB9, 8'h88, 8'h00, 8'h30, 8'h13, 8'hB9, 8'hBD, 8'h00, 8'hD0, 8'h0E, 8'hA9, 8'h00, 8'h95, 8'h31, 8'hB9,
			8'h9A, 8'h00, 8'h38, 8'hE9, 8'h04, 8'hD5, 8'h9A, 8'hB0, 8'h04, 8'hA9, 8'h40, 8'h95, 8'h31, 8'hB5, 8'h91, 8'hD9,
			8'h91, 8'h00, 8'hB0, 8'h07, 8'hB5, 8'h31, 8'h09, 8'h01, 8'h95, 8'h31, 8'h60, 8'hB5, 8'h31, 8'h09, 8'h02, 8'h95,
			8'h31, 8'h60, 8'h1F, 8'h0F, 8'h07, 8'h20, 8'h10, 8'h08, 8'hA2, 8'h00, 8'hA9, 8'h01, 8'h8D, 8'h16, 8'h40, 8'hA9,
			8'h00, 8'h8D, 8'h16, 8'h40, 8'hA0, 8'h07, 8'hBD, 8'h16, 8'h40, 8'h85, 8'h12, 8'h4A, 8'h05, 8'h12, 8'h4A, 8'h3E,
			8'h1C, 8'h06, 8'h88, 8'h10, 8'hF1, 8'hBC, 8'h1E, 8'h06, 8'hBD, 8'h1C, 8'h06, 8'h9D, 8'h1E, 8'h06, 8'h98, 8'h5D,
			8'h1C, 8'h06, 8'h3D, 8'h1C, 8'h06, 8'h60, 8'hB5, 8'h88, 8'hD0, 8'h09, 8'hA9, 8'h00, 8'h9D, 8'h24, 8'h04, 8'h9D,
			8'h2D, 8'h04, 8'h60, 8'hC9, 8'h02, 8'hF0, 8'h41, 8'hE0, 8'h02, 8'h90, 8'h3D, 8'hB5, 8'h7F, 8'hC9, 8'h02, 8'hB0,
			8'hE9, 8'hBD, 8'h24, 8'h04, 8'h85, 8'h12, 8'hBD, 8'h2D, 8'h04, 8'h85, 8'h13, 8'h20, 8'hA6, 8'hF1, 8'hBD, 8'h63,
			8'h04, 8'h18, 8'h65, 8'h12, 8'h9D, 8'h63, 8'h04, 8'h85, 8'h12, 8'hBD, 8'h6C, 8'h04, 8'h65, 8'h13, 8'h9D, 8'h6C,
			8'h04, 8'h85, 8'h13, 8'h20, 8'hA6, 8'hF1, 8'hBD, 8'h24, 8'h04, 8'h38, 8'hE5, 8'h12, 8'h9D, 8'h24, 8'h04, 8'hBD,
			8'h2D, 8'h04, 8'hE5, 8'h13, 8'h9D, 8'h2D, 8'h04, 8'h60, 8'hB5, 8'h7F, 8'hC9, 8'h06, 8'h90, 8'h01, 8'h60, 8'hB5,
			8'h7F, 8'hC9, 8'h04, 8'hD0, 8'h1C, 8'hB5, 8'h31, 8'h29, 8'h02, 8'hF0, 8'h07, 8'hBD, 8'h48, 8'h04, 8'hF0, 8'h11,
			8'hD0, 8'h0B, 8'hB5, 8'h31, 8'h29, 8'h01, 8'hF0, 8'h09, 8'hBD, 8'h48, 8'h04, 8'hD0, 8'h04, 8'hA9, 8'h05, 8'h95,
			8'h7F, 8'hB5, 8'h7F, 8'hC9, 8'h02, 8'hD0, 8'h1B, 8'hB5, 8'h31, 8'h29, 8'h02, 8'hF0, 8'h04, 8'hA9, 8'h00, 8'hF0,
			8'h08, 8'hB5, 8'h31, 8'h29, 8'h01, 8'hF0, 8'h07, 8'hA9, 8'h01, 8'hDD, 8'h48, 8'h04, 8'hF0, 8'h04, 8'hA9, 8'h04,
			8'h95, 8'h7F, 8'hB5, 8'h7F, 8'hC9, 8'h04, 8'h90, 8'h1C, 8'hB5, 8'h31, 8'h29, 8'h02, 8'hF0, 8'h07, 8'hBD, 8'h48,
			8'h04, 8'hD0, 8'h11, 8'hF0, 8'h0B, 8'hB5, 8'h31, 8'h29, 8'h01, 8'hF0, 8'h09, 8'hBD, 8'h48, 8'h04, 8'hF0, 8'h04,
			8'hA9, 8'h02, 8'h95, 8'h7F, 8'hB5, 8'h7F, 8'hC9, 8'h03, 8'hD0, 8'h0A, 8'hB5, 8'h31, 8'h29, 8'h03, 8'hF0, 8'h04,
			8'hA9, 8'h02, 8'h95, 8'h7F, 8'hB5, 8'h7F, 8'hC9, 8'h04, 8'hB0, 8'h15, 8'hB5, 8'h31, 8'h29, 8'h02, 8'hF0, 8'h04,
			8'hA9, 8'h00, 8'hF0, 8'h08, 8'hB5, 8'h31, 8'h29, 8'h01, 8'hF0, 8'h05, 8'hA9, 8'h01, 8'h9D, 8'h48, 8'h04, 8'hB5,
			8'h7F, 8'hC9, 8'h04, 8'h90, 8'h33, 8'hBD, 8'h36, 8'h04, 8'hC9, 8'h01, 8'hD0, 8'h2C, 8'hBC, 8'h51, 8'h04, 8'hBD,
			8'h48, 8'h04, 8'hF0, 8'h12, 8'hBD, 8'h24, 8'h04, 8'h38, 8'hF9, 8'h25, 8'hE6, 8'h9D, 8'h24, 8'h04, 8'hBD, 8'h2D,
			8'h04, 8'hE9, 8'h00, 8'h4C, 8'h01, 8'hE9, 8'hBD, 8'h24, 8'h04, 8'h18, 8'h79, 8'h25, 8'hE6, 8'h9D, 8'h24, 8'h04,
			8'hBD, 8'h2D, 8'h04, 8'h69, 8'h00, 8'h4C, 8'h01, 8'hE9, 8'hB5, 8'h7F, 8'hF0, 8'h0B, 8'hC9, 8'h02, 8'hF0, 8'h47,
			8'hC9, 8'h03, 8'hF0, 8'h03, 8'h4C, 8'h51, 8'hE9, 8'hBD, 8'h36, 8'h04, 8'hC9, 8'h01, 8'hF0, 8'h03, 8'h4C, 8'h51,
			8'hE9, 8'hBC, 8'h51, 8'h04, 8'hB5, 8'h31, 8'h29, 8'h02, 8'hF0, 8'h12, 8'hBD, 8'h24, 8'h04, 8'h38, 8'hF9, 8'h19,
			8'hE6, 8'h9D, 8'h24, 8'h04, 8'hBD, 8'h2D, 8'h04, 8'hE9, 8'h00, 8'h4C, 8'h01, 8'hE9, 8'hB5, 8'h31, 8'h29, 8'h01,
			8'hF0, 8'h5F, 8'hBD, 8'h24, 8'h04, 8'h18, 8'h79, 8'h19, 8'hE6, 8'h9D, 8'h24, 8'h04, 8'hBD, 8'h2D, 8'h04, 8'h69,
			8'h00, 8'h9D, 8'h2D, 8'h04, 8'h4C, 8'h51, 8'hE9, 8'hBD, 8'h36, 8'h04, 8'hC9, 8'h01, 8'hD0, 8'h43, 8'hBC, 8'h51,
			8'h04, 8'hB5, 8'h31, 8'h29, 8'h02, 8'hF0, 8'h12, 8'hBD, 8'h24, 8'h04, 8'h38, 8'hF9, 8'h25, 8'hE6, 8'h9D, 8'h24,
			8'h04, 8'hBD, 8'h2D, 8'h04, 8'hE9, 8'h00, 8'h4C, 8'h3E, 8'hE9, 8'hB5, 8'h31, 8'h29, 8'h01, 8'hF0, 8'h22, 8'hBD,
			8'h24, 8'h04, 8'h18, 8'h79, 8'h25, 8'hE6, 8'h9D, 8'h24, 8'h04, 8'hBD, 8'h2D, 8'h04, 8'h69, 8'h00, 8'h9D, 8'h2D,
			8'h04, 8'hB5, 8'h31, 8'h29, 8'h03, 8'hF0, 8'h0A, 8'hE0, 8'h02, 8'hB0, 8'h06, 8'hA5, 8'hF0, 8'h09, 8'h08, 8'h85,
			8'hF0, 8'hB5, 8'h7F, 8'hC9, 8'h04, 8'h90, 8'h2B, 8'hBD, 8'h48, 8'h04, 8'hD0, 8'h07, 8'hBD, 8'h2D, 8'h04, 8'h30,
			8'h21, 8'h10, 8'h05, 8'hBD, 8'h2D, 8'h04, 8'h10, 8'h1A, 8'hB5, 8'h7F, 8'hC9, 8'h05, 8'hD0, 8'h08, 8'hBD, 8'h48,
			8'h04, 8'h49, 8'h01, 8'h9D, 8'h48, 8'h04, 8'hA9, 8'h03, 8'h95, 8'h7F, 8'hA9, 8'h00, 8'h9D, 8'h24, 8'h04, 8'h9D,
			8'h2D, 8'h04, 8'h60, 8'hA5, 8'hCB, 8'hD0, 8'h2F, 8'hB5, 8'hBD, 8'hF0, 8'h0F, 8'hAD, 8'h88, 8'h04, 8'hF0, 8'h0A,
			8'h38, 8'hF5, 8'h91, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h05, 8'h90, 8'h1C, 8'hE0, 8'h02, 8'h90, 8'h06, 8'hB5, 8'h88,
			8'hC9, 8'h02, 8'hD0, 8'h4E, 8'hB5, 8'h7F, 8'hC9, 8'h02, 8'h90, 8'h48, 8'hC9, 8'h06, 8'hB0, 8'h44, 8'hA9, 8'h01,
			8'h95, 8'h7F, 8'h9D, 8'h5A, 8'h04, 8'h60, 8'hA9, 8'h00, 8'h9D, 8'h12, 8'h04, 8'h9D, 8'h1B, 8'h04, 8'h9D, 8'h09,
			8'h04, 8'h85, 8'hCB, 8'hE0, 8'h02, 8'h90, 8'h36, 8'hB5, 8'h88, 8'hC9, 8'h02, 8'hF0, 8'h26, 8'hC9, 8'h01, 8'hD0,
			8'h21, 8'hB5, 8'h7F, 8'hC9, 8'h02, 8'hB0, 8'h1B, 8'hA9, 8'h02, 8'h95, 8'h7F, 8'hA5, 8'hC6, 8'h9D, 8'h3F, 8'h04,
			8'hA9, 8'h00, 8'h9D, 8'h24, 8'h04, 8'h9D, 8'h2D, 8'h04, 8'h9D, 8'h63, 8'h04, 8'h9D, 8'h6C, 8'h04, 8'hA9, 8'h40,
			8'h85, 8'hF1, 8'h60, 8'hA9, 8'h00, 8'h95, 8'h7F, 8'hA9, 8'h01, 8'h9D, 8'h5A, 8'h04, 8'h60, 8'hB5, 8'h7F, 8'hC9,
			8'h01, 8'hD0, 8'h14, 8'hC9, 8'h06, 8'hB0, 8'h10, 8'hBD, 8'h24, 8'h04, 8'h1D, 8'h2D, 8'h04, 8'hD0, 8'h04, 8'hA9,
			8'h03, 8'hD0, 8'h02, 8'hA9, 8'h02, 8'h95, 8'h7F, 8'h60, 8'hE0, 8'h02, 8'hB0, 8'h10, 8'hB5, 8'hBD, 8'hD0, 8'h24,
			8'hB5, 8'h7F, 8'hC9, 8'h01, 8'hF0, 8'h18, 8'hC9, 8'h03, 8'hD0, 8'h1A, 8'hF0, 8'h12, 8'hB5, 8'h7F, 8'hC9, 8'h01,
			8'hF0, 8'h0C, 8'hC9, 8'h03, 8'h90, 8'h0E, 8'hA5, 8'h19, 8'h29, 8'h03, 8'hD0, 8'h0B, 8'hF0, 8'h06, 8'hA5, 8'h19,
			8'h29, 8'h07, 8'hD0, 8'h03, 8'hFE, 8'h36, 8'h04, 8'hBD, 8'h36, 8'h04, 8'h29, 8'h03, 8'h9D, 8'h36, 8'h04, 8'hD0,
			8'h06, 8'hB5, 8'h7F, 8'hD0, 8'h02, 8'hF6, 8'h7F, 8'h60, 8'hBD, 8'h75, 8'h04, 8'hF0, 8'h03, 8'hDE, 8'h75, 8'h04,
			8'hE0, 8'h02, 8'hB0, 8'h28, 8'hB5, 8'hC1, 8'hF0, 8'h24, 8'hA5, 8'h19, 8'h4A, 8'h90, 8'h1E, 8'hFE, 8'h36, 8'h04,
			8'hBD, 8'h36, 8'h04, 8'h29, 8'h03, 8'h9D, 8'h36, 8'h04, 8'hA9, 8'h01, 8'h95, 8'h7F, 8'hDE, 8'h5A, 8'h04, 8'hD0,
			8'h0A, 8'hA9, 8'h00, 8'h95, 8'hC1, 8'h95, 8'h7F, 8'hA9, 8'h20, 8'h85, 8'hF0, 8'h60, 8'hBD, 8'h12, 8'h04, 8'h18,
			8'hBC, 8'h51, 8'h04, 8'h79, 8'h01, 8'hE6, 8'h9D, 8'h12, 8'h04, 8'h90, 8'h03, 8'hFE, 8'h1B, 8'h04, 8'hBD, 8'h1B,
			8'h04, 8'h30, 8'h1E, 8'hD9, 8'h6D, 8'hE6, 8'h90, 8'h34, 8'hD0, 8'h08, 8'hBD, 8'h12, 8'h04, 8'hD9, 8'h61, 8'hE6,
			8'h90, 8'h2A, 8'hB9, 8'h61, 8'hE6, 8'h9D, 8'h12, 8'h04, 8'hB9, 8'h6D, 8'hE6, 8'h9D, 8'h1B, 8'h04, 8'h4C, 8'hDC,
			8'hEA, 8'hD9, 8'h85, 8'hE6, 8'h90, 8'h0A, 8'hD0, 8'h14, 8'hBD, 8'h12, 8'h04, 8'hD9, 8'h79, 8'hE6, 8'hB0, 8'h0C,
			8'hB9, 8'h79, 8'hE6, 8'h9D, 8'h12, 8'h04, 8'hB9, 8'h85, 8'hE6, 8'h9D, 8'h1B, 8'h04, 8'h20, 8'hA0, 8'hEB, 8'hC9,
			8'hF8, 8'hB0, 8'h2A, 8'hC9, 8'hE8, 8'h90, 8'h26, 8'hA9, 8'hFF, 8'h95, 8'h88, 8'hA9, 8'h04, 8'h85, 8'hBB, 8'hB5,
			8'h91, 8'h85, 8'hBC, 8'hE0, 8'h02, 8'h90, 8'h0E, 8'hA9, 8'h80, 8'h95, 8'h88, 8'hA9, 8'h00, 8'h95, 8'h7F, 8'hA9,
			8'h01, 8'h85, 8'hF3, 8'hD0, 8'h08, 8'hA5, 8'hC8, 8'hD0, 8'h04, 8'hA9, 8'h40, 8'h85, 8'hF0, 8'hBD, 8'h2D, 8'h04,
			8'h30, 8'h1E, 8'hD9, 8'h3D, 8'hE6, 8'h90, 8'h34, 8'hD0, 8'h08, 8'hBD, 8'h24, 8'h04, 8'hD9, 8'h31, 8'hE6, 8'h90,
			8'h2A, 8'hB9, 8'h31, 8'hE6, 8'h9D, 8'h24, 8'h04, 8'hB9, 8'h3D, 8'hE6, 8'h9D, 8'h2D, 8'h04, 8'h4C, 8'h4B, 8'hEB,
			8'hD9, 8'h55, 8'hE6, 8'h90, 8'h0A, 8'hD0, 8'h14, 8'hBD, 8'h24, 8'h04, 8'hD9, 8'h49, 8'hE6, 8'hB0, 8'h0C, 8'hB9,
			8'h49, 8'hE6, 8'h9D, 8'h24, 8'h04, 8'hB9, 8'h55, 8'hE6, 8'h9D, 8'h2D, 8'h04, 8'h20, 8'h8E, 8'hEB, 8'hA5, 8'h16,
			8'hF0, 8'h10, 8'hB5, 8'h91, 8'hC9, 8'h10, 8'hB0, 8'h02, 8'hA9, 8'h10, 8'hC9, 8'hE0, 8'h90, 8'h02, 8'hA9, 8'hE0,
			8'h95, 8'h91, 8'hA5, 8'hC8, 8'hF0, 8'h27, 8'hB5, 8'h88, 8'hD0, 8'h23, 8'hB5, 8'h9A, 8'hC9, 8'hC8, 8'h90, 8'h1D,
			8'hA9, 8'hC7, 8'h95, 8'h9A, 8'hBD, 8'h51, 8'h04, 8'hC9, 8'h0B, 8'hD0, 8'h09, 8'hDE, 8'h51, 8'h04, 8'h20, 8'h07,
			8'hF1, 8'h4C, 8'h8C, 8'hF1, 8'hA9, 8'h02, 8'h95, 8'h88, 8'hA9, 8'h03, 8'h9D, 8'h51, 8'h04, 8'h60, 8'hBD, 8'h00,
			8'h04, 8'h18, 8'h7D, 8'h24, 8'h04, 8'h9D, 8'h00, 8'h04, 8'hB5, 8'h91, 8'h7D, 8'h2D, 8'h04, 8'h95, 8'h91, 8'h60,
			8'hBD, 8'h09, 8'h04, 8'h18, 8'h7D, 8'h12, 8'h04, 8'h9D, 8'h09, 8'h04, 8'hB5, 8'h9A, 8'h7D, 8'h1B, 8'h04, 8'h95,
			8'h9A, 8'h60, 8'h20, 8'hB4, 8'hF0, 8'h20, 8'h8E, 8'hEB, 8'h4C, 8'hB4, 8'hF0, 8'h20, 8'hB4, 8'hF0, 8'h20, 8'hA0,
			8'hEB, 8'h4C, 8'hB4, 8'hF0, 8'hE0, 8'h02, 8'hB0, 8'h1B, 8'hB5, 8'h88, 8'hD0, 8'h0A, 8'hBD, 8'h36, 8'h04, 8'hD0,
			8'h05, 8'hA9, 8'h00, 8'h95, 8'h7F, 8'h60, 8'hB5, 8'h7F, 8'hC9, 8'h06, 8'h90, 8'h5C, 8'hA9, 8'h01, 8'h95, 8'h7F,
			8'hD6, 8'h88, 8'h60, 8'hB5, 8'h88, 8'hC9, 8'h02, 8'hF0, 8'h4F, 8'hBD, 8'h36, 8'h04, 8'hD0, 8'h0F, 8'hB5, 8'h88,
			8'hD0, 8'h05, 8'hA9, 8'h00, 8'h95, 8'h7F, 8'h60, 8'hB5, 8'h7F, 8'hD0, 8'h03, 8'hF6, 8'h7F, 8'h60, 8'hC9, 8'h02,
			8'h90, 8'hFB, 8'hDE, 8'h5A, 8'h04, 8'hD0, 8'h30, 8'hA5, 8'hC7, 8'h9D, 8'h5A, 8'h04, 8'hF6, 8'h7F, 8'hB5, 8'h7F,
			8'hC9, 8'h07, 8'h90, 8'h23, 8'hA9, 8'h02, 8'h95, 8'h88, 8'hA9, 8'h00, 8'h95, 8'h7F, 8'hBC, 8'h51, 8'h04, 8'hB9,
			8'hAE, 8'hEC, 8'hBC, 8'h7E, 8'h04, 8'hD0, 8'h08, 8'hDE, 8'h7E, 8'h04, 8'hBD, 8'h51, 8'h04, 8'h29, 8'h03, 8'h9D,
			8'h51, 8'h04, 8'hA9, 8'hFE, 8'h9D, 8'h1B, 8'h04, 8'h60, 8'h20, 8'hE9, 8'hE6, 8'hB5, 8'h31, 8'h29, 8'hC3, 8'hF0,
			8'h08, 8'hE0, 8'h02, 8'hB0, 8'h04, 8'hA9, 8'h00, 8'h95, 8'hBD, 8'hB5, 8'h31, 8'h29, 8'h40, 8'hD0, 8'h12, 8'hB5,
			8'h31, 8'h29, 8'h80, 8'hD0, 8'h07, 8'hA9, 8'h00, 8'h9D, 8'h20, 8'h06, 8'hF0, 8'h51, 8'hBD, 8'h20, 8'h06, 8'hD0,
			8'h4C, 8'hB5, 8'h7F, 8'hC9, 8'h02, 8'h90, 8'h0E, 8'hD6, 8'h9A, 8'hD6, 8'h9A, 8'hA9, 8'h00, 8'h9D, 8'h12, 8'h04,
			8'h9D, 8'h1B, 8'h04, 8'hF0, 8'h09, 8'hC9, 8'h01, 8'hF0, 8'h05, 8'hBD, 8'h36, 8'h04, 8'hD0, 8'h2F, 8'hA9, 8'h00,
			8'h95, 8'h7F, 8'hA9, 8'h01, 8'h9D, 8'h36, 8'h04, 8'hA9, 8'h01, 8'h9D, 8'h20, 8'h06, 8'hA0, 8'h00, 8'hE0, 8'h02,
			8'h90, 8'h01, 8'hC8, 8'hB9, 8'hF0, 8'h00, 8'h09, 8'h10, 8'h99, 8'hF0, 8'h00, 8'hBD, 8'h12, 8'h04, 8'h38, 8'hBC,
			8'h51, 8'h04, 8'hF9, 8'h0D, 8'hE6, 8'h9D, 8'h12, 8'h04, 8'hB0, 8'h03, 8'hDE, 8'h1B, 8'h04, 8'h60, 8'h01, 8'h02,
			8'h02, 8'h03, 8'h01, 8'h02, 8'h02, 8'h03, 8'h01, 8'h02, 8'h02, 8'h03, 8'hB5, 8'h7F, 8'hD0, 8'h69, 8'h20, 8'hB1,
			8'hE7, 8'h20, 8'h8E, 8'hEB, 8'hBD, 8'h09, 8'h04, 8'h38, 8'hE9, 8'h60, 8'h9D, 8'h09, 8'h04, 8'hB5, 8'h9A, 8'hE9,
			8'h00, 8'h95, 8'h9A, 8'hC9, 8'hF1, 8'h90, 8'h04, 8'hA9, 8'hFF, 8'h95, 8'h88, 8'h8A, 8'h48, 8'hA0, 8'h01, 8'hB9,
			8'h88, 8'h00, 8'hF0, 8'h3E, 8'h30, 8'h3C, 8'hB5, 8'h9A, 8'h38, 8'hF9, 8'h9A, 8'h00, 8'h20, 8'h8E, 8'hF0, 8'hC9,
			8'h18, 8'hB0, 8'h2F, 8'hB5, 8'h91, 8'h38, 8'hF9, 8'h91, 8'h00, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h10, 8'hB0, 8'h22,
			8'hA9, 8'hFF, 8'h95, 8'h7F, 8'hA9, 8'h03, 8'h9D, 8'h5A, 8'h04, 8'hA9, 8'h78, 8'h85, 8'hC5, 8'hA9, 8'h02, 8'h85,
			8'hF0, 8'hA9, 8'h32, 8'h84, 8'h3E, 8'h20, 8'hDE, 8'hD6, 8'hA9, 8'h01, 8'hA6, 8'h3E, 8'h20, 8'h71, 8'hD8, 8'h68,
			8'hAA, 8'h60, 8'h88, 8'h10, 8'hBA, 8'h68, 8'hAA, 8'h60, 8'hB4, 8'h88, 8'h88, 8'h10, 8'h01, 8'h60, 8'hB5, 8'h9A,
			8'hC9, 8'hF9, 8'h90, 8'h0C, 8'hBD, 8'h1B, 8'h04, 8'h10, 8'hF4, 8'hA9, 8'h00, 8'h85, 8'hCC, 8'h4C, 8'hE1, 8'hED,
			8'hA4, 8'hCD, 8'h30, 8'hE3, 8'hA9, 8'h00, 8'h85, 8'hCC, 8'hB1, 8'h27, 8'h38, 8'hE9, 8'h18, 8'hD5, 8'h9A, 8'hB0,
			8'h65, 8'h69, 8'h03, 8'hD5, 8'h9A, 8'h90, 8'h04, 8'hA9, 8'h01, 8'hD0, 8'h0E, 8'hB1, 8'h29, 8'hD5, 8'h9A, 8'h90,
			8'h55, 8'hE9, 8'h03, 8'hD5, 8'h9A, 8'hB0, 8'h22, 8'hA9, 8'h02, 8'h85, 8'hCC, 8'hB1, 8'h23, 8'hC9, 8'h10, 8'hF0,
			8'h07, 8'h38, 8'hE9, 8'h0C, 8'hD5, 8'h91, 8'hB0, 8'h0D, 8'hB1, 8'h25, 8'hC9, 8'hFF, 8'hF0, 8'h0B, 8'h38, 8'hE9,
			8'h04, 8'hD5, 8'h91, 8'hB0, 8'h04, 8'hA9, 8'h00, 8'h85, 8'hCC, 8'hB1, 8'h23, 8'h38, 8'hE9, 8'h10, 8'hF0, 8'h10,
			8'hD5, 8'h91, 8'hB0, 8'h22, 8'h69, 8'h04, 8'hD5, 8'h91, 8'h90, 8'h06, 8'hA5, 8'hCC, 8'h09, 8'h04, 8'hD0, 8'h14,
			8'hB1, 8'h25, 8'hC9, 8'hFF, 8'hF0, 8'h10, 8'hD5, 8'h91, 8'h90, 8'h0C, 8'hE9, 8'h04, 8'hD5, 8'h91, 8'hB0, 8'h06,
			8'hA5, 8'hCC, 8'h09, 8'h08, 8'h85, 8'hCC, 8'hA5, 8'hCC, 8'hD0, 8'h07, 8'h88, 8'h30, 8'h03, 8'h4C, 8'h44, 8'hED,
			8'h60, 8'h46, 8'hCC, 8'h90, 8'h11, 8'hBD, 8'h1B, 8'h04, 8'h30, 8'h0C, 8'hB1, 8'h27, 8'hE9, 8'h18, 8'h95, 8'h9A,
			8'hF6, 8'h9A, 8'hA9, 8'h01, 8'h85, 8'hCB, 8'h46, 8'hCC, 8'h90, 8'h1A, 8'hBD, 8'h1B, 8'h04, 8'h10, 8'h15, 8'hB1,
			8'h29, 8'h95, 8'h9A, 8'h20, 8'h07, 8'hF1, 8'h20, 8'h8C, 8'hF1, 8'hE0, 8'h02, 8'hB0, 8'h03, 8'h20, 8'h33, 8'hCC,
			8'hA5, 8'hCB, 8'hD0, 8'h30, 8'h46, 8'hCC, 8'h90, 8'h07, 8'hBD, 8'h2D, 8'h04, 8'h30, 8'h02, 8'h10, 8'h09, 8'h46,
			8'hCC, 8'h90, 8'h21, 8'hBD, 8'h2D, 8'h04, 8'h10, 8'h1C, 8'h20, 8'hDE, 8'hF0, 8'h20, 8'h72, 8'hF1, 8'hBD, 8'h2D,
			8'h04, 8'h1D, 8'h24, 8'h04, 8'hF0, 8'h0E, 8'hBD, 8'h48, 8'h04, 8'h49, 8'h01, 8'h9D, 8'h48, 8'h04, 8'hA5, 8'hF1,
			8'h09, 8'h02, 8'h85, 8'hF1, 8'h60, 8'hA2, 8'h07, 8'h86, 8'h12, 8'hA4, 8'h12, 8'h88, 8'h10, 8'h03, 8'h4C, 8'h2A,
			8'hEF, 8'hB5, 8'h88, 8'h30, 8'hF9, 8'hF0, 8'hF7, 8'hB9, 8'h88, 8'h00, 8'h30, 8'hF2, 8'hF0, 8'hF0, 8'hA9, 8'h00,
			8'h85, 8'hCC, 8'hB9, 8'h9A, 8'h00, 8'h38, 8'hF5, 8'h9A, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h18, 8'hB0, 8'h71, 8'hB5,
			8'h9A, 8'h18, 8'h69, 8'h18, 8'h85, 8'h12, 8'hB9, 8'h9A, 8'h00, 8'h18, 8'h69, 8'h07, 8'h38, 8'hE5, 8'h12, 8'h20,
			8'h8E, 8'hF0, 8'hC9, 8'h04, 8'hB0, 8'h04, 8'hA9, 8'h01, 8'hD0, 8'h12, 8'hB9, 8'h9A, 8'h00, 8'h18, 8'h69, 8'h11,
			8'h38, 8'hF5, 8'h9A, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h04, 8'hB0, 8'h15, 8'hA9, 8'h02, 8'h85, 8'hCC, 8'hB9, 8'h91,
			8'h00, 8'h38, 8'hF5, 8'h91, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h10, 8'h90, 8'h04, 8'hA9, 8'h00, 8'h85, 8'hCC, 8'hB5,
			8'h91, 8'h18, 8'h69, 8'h10, 8'h85, 8'h12, 8'hB9, 8'h91, 8'h00, 8'h18, 8'h69, 8'h07, 8'h38, 8'hE5, 8'h12, 8'h20,
			8'h8E, 8'hF0, 8'hC9, 8'h04, 8'hB0, 8'h04, 8'hA9, 8'h04, 8'hD0, 8'h12, 8'hB9, 8'h91, 8'h00, 8'h18, 8'h69, 8'h09,
			8'h38, 8'hF5, 8'h91, 8'h20, 8'h8E, 8'hF0, 8'hC9, 8'h04, 8'hB0, 8'h06, 8'hA9, 8'h08, 8'h05, 8'hCC, 8'h85, 8'hCC,
			8'hA9, 8'h00, 8'h85, 8'h4B, 8'h46, 8'hCC, 8'h90, 8'h05, 8'h20, 8'hA6, 8'hF0, 8'h30, 8'h09, 8'h46, 8'hCC, 8'h90,
			8'h20, 8'h20, 8'hA6, 8'hF0, 8'h30, 8'h1B, 8'h20, 8'hBD, 8'hF0, 8'hB0, 8'h12, 8'h20, 8'h07, 8'hF1, 8'h20, 8'h8C,
			8'hF1, 8'h20, 8'hB4, 8'hF0, 8'h20, 8'h07, 8'hF1, 8'h20, 8'h8C, 8'hF1, 8'h20, 8'hB4, 8'hF0, 8'hA9, 8'h01, 8'h85,
			8'h4B, 8'h46, 8'hCC, 8'h90, 8'h05, 8'h20, 8'h98, 8'hF0, 8'h30, 8'h09, 8'h46, 8'hCC, 8'h90, 8'h20, 8'h20, 8'h98,
			8'hF0, 8'h30, 8'h1B, 8'h20, 8'hBD, 8'hF0, 8'hB0, 8'h12, 8'h20, 8'hDE, 8'hF0, 8'h20, 8'h72, 8'hF1, 8'h20, 8'hB4,
			8'hF0, 8'h20, 8'hDE, 8'hF0, 8'h20, 8'h72, 8'hF1, 8'h20, 8'hB4, 8'hF0, 8'hA9, 8'h01, 8'h85, 8'h4B, 8'h20, 8'h37,
			8'hEF, 8'h20, 8'hB4, 8'hF0, 8'h20, 8'h37, 8'hEF, 8'h20, 8'hB4, 8'hF0, 8'h88, 8'h30, 8'h03, 8'h4C, 8'h31, 8'hEE,
			8'hCA, 8'h30, 8'h03, 8'h4C, 8'h27, 8'hEE, 8'h60, 8'hE0, 8'h02, 8'h90, 8'h07, 8'hC0, 8'h02, 8'h90, 8'h03, 8'h4C,
			8'h43, 8'hF0, 8'hA9, 8'h00, 8'h8D, 8'h87, 8'h04, 8'hBD, 8'h75, 8'h04, 8'hF0, 8'h03, 8'h4C, 8'h43, 8'hF0, 8'hA5,
			8'h4B, 8'hD0, 8'h03, 8'h4C, 8'h43, 8'hF0, 8'hE0, 8'h02, 8'hB0, 8'h07, 8'hB5, 8'hBD, 8'hF0, 8'h14, 8'h4C, 8'h43,
			8'hF0, 8'hB5, 8'h88, 8'hC9, 8'h01, 8'hD0, 8'h0B, 8'hB5, 8'h7F, 8'hC9, 8'h02, 8'hB0, 8'h12, 8'hA9, 8'h01, 8'h8D,
			8'h87, 8'h04, 8'hB9, 8'h9A, 8'h00, 8'h18, 8'h69, 8'h04, 8'hD5, 8'h9A, 8'h90, 8'h03, 8'h4C, 8'h43, 8'hF0, 8'hA9,
			8'h14, 8'h9D, 8'h75, 8'h04, 8'hA9, 8'h00, 8'h9D, 8'h36, 8'h04, 8'hC0, 8'h02, 8'h90, 8'h0A, 8'hB9, 8'h88, 8'h00,
			8'hC9, 8'h02, 8'hF0, 8'h03, 8'h4C, 8'h43, 8'hF0, 8'hA5, 8'hF0, 8'h09, 8'h02, 8'h85, 8'hF0, 8'hB5, 8'h88, 8'hC9,
			8'h02, 8'hD0, 8'h1D, 8'hE0, 8'h02, 8'hB0, 8'h19, 8'h84, 8'h12, 8'hB4, 8'h7F, 8'hB9, 8'h53, 8'hF0, 8'hA4, 8'h12,
			8'h48, 8'h68, 8'hD0, 8'h03, 8'h4C, 8'h43, 8'hF0, 8'h95, 8'h7F, 8'hA9, 8'h00, 8'h9D, 8'h36, 8'h04, 8'hF0, 8'h2A,
			8'hD6, 8'h88, 8'hD0, 8'h0A, 8'hA9, 8'hFF, 8'h9D, 8'h1B, 8'h04, 8'hA9, 8'h00, 8'h9D, 8'h12, 8'h04, 8'hA9, 8'h00,
			8'h95, 8'h7F, 8'h9D, 8'h24, 8'h04, 8'h9D, 8'h2D, 8'h04, 8'hB5, 8'h91, 8'h30, 8'h04, 8'hA9, 8'hFF, 8'hD0, 8'h02,
			8'hA9, 8'h00, 8'h9D, 8'h6C, 8'h04, 8'hA9, 8'h80, 8'h9D, 8'h63, 8'h04, 8'h84, 8'h12, 8'hBC, 8'h51, 8'h04, 8'hB9,
			8'h5E, 8'hF0, 8'h9D, 8'h51, 8'h04, 8'hA9, 8'h01, 8'h9D, 8'h7E, 8'h04, 8'hA4, 8'h12, 8'hC0, 8'h02, 8'hB0, 8'h43,
			8'hBD, 8'h51, 8'h04, 8'hC9, 8'h07, 8'hF0, 8'h0A, 8'hC9, 8'h08, 8'h90, 8'h06, 8'hA5, 8'hF1, 8'h09, 8'h80, 8'h85,
			8'hF1, 8'hBC, 8'h51, 8'h04, 8'hB9, 8'h6A, 8'hF0, 8'h85, 8'h13, 8'hAD, 8'h87, 8'h04, 8'hF0, 8'h05, 8'hB9, 8'h76,
			8'hF0, 8'h85, 8'h13, 8'hB9, 8'h82, 8'hF0, 8'h18, 8'h6D, 8'h87, 8'h04, 8'h85, 8'h14, 8'hA5, 8'h12, 8'h85, 8'h3E,
			8'h48, 8'h8A, 8'h48, 8'hA5, 8'h13, 8'h48, 8'hA5, 8'h14, 8'h20, 8'h71, 8'hD8, 8'h68, 8'h20, 8'hDE, 8'hD6, 8'h68,
			8'hAA, 8'h68, 8'hA8, 8'hBD, 8'h51, 8'h04, 8'hC9, 8'h0B, 8'hD0, 8'h08, 8'hA5, 8'hC8, 8'hD0, 8'h04, 8'hA9, 8'h20,
			8'h85, 8'hF0, 8'h60, 8'h06, 8'h06, 8'h07, 8'h08, 8'h09, 8'h0A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h05,
			8'h06, 8'h07, 8'h08, 8'h09, 8'h0A, 8'h0B, 8'h08, 8'h09, 8'h0A, 8'h0B, 8'h00, 8'h00, 8'h00, 8'h00, 8'h32, 8'h4B,
			8'h64, 8'h64, 8'h4B, 8'h64, 8'h96, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h32, 8'h4B, 8'h64, 8'h64, 8'h64, 8'h96,
			8'hC8, 8'h64, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h02, 8'h03, 8'h03, 8'h02, 8'h03, 8'h04, 8'h03, 8'h48, 8'h68,
			8'h10, 8'h05, 8'h49, 8'hFF, 8'h18, 8'h69, 8'h01, 8'h60, 8'hB9, 8'h24, 8'h04, 8'h38, 8'hFD, 8'h24, 8'h04, 8'hB9,
			8'h2D, 8'h04, 8'hFD, 8'h2D, 8'h04, 8'h60, 8'hB9, 8'h12, 8'h04, 8'h38, 8'hFD, 8'h12, 8'h04, 8'hB9, 8'h1B, 8'h04,
			8'hFD, 8'h1B, 8'h04, 8'h60, 8'h86, 8'h12, 8'h84, 8'h13, 8'hA6, 8'h13, 8'hA4, 8'h12, 8'h60, 8'hE0, 8'h02, 8'h90,
			8'h1C, 8'hB5, 8'h7F, 8'hC9, 8'h02, 8'h90, 8'h16, 8'hA9, 8'h01, 8'hD5, 8'h88, 8'hB0, 8'h10, 8'hC0, 8'h02, 8'h90,
			8'h0C, 8'hB9, 8'h7F, 8'h00, 8'hC9, 8'h02, 8'h90, 8'h05, 8'hA9, 8'h01, 8'hD9, 8'h88, 8'h00, 8'h60, 8'hA9, 8'h00,
			8'h38, 8'hFD, 8'h24, 8'h04, 8'h9D, 8'h24, 8'h04, 8'hA9, 8'h00, 8'hFD, 8'h2D, 8'h04, 8'h9D, 8'h2D, 8'h04, 8'hA9,
			8'h00, 8'h38, 8'hFD, 8'h63, 8'h04, 8'h9D, 8'h63, 8'h04, 8'hA9, 8'h00, 8'hFD, 8'h6C, 8'h04, 8'h9D, 8'h6C, 8'h04,
			8'hB5, 8'h31, 8'h29, 8'h40, 8'h95, 8'h31, 8'h60, 8'hA9, 8'h00, 8'h38, 8'hFD, 8'h12, 8'h04, 8'h9D, 8'h12, 8'h04,
			8'hA9, 8'h00, 8'hFD, 8'h1B, 8'h04, 8'h9D, 8'h1B, 8'h04, 8'h60, 8'h85, 8'h2D, 8'hA5, 8'h2C, 8'h10, 8'h24, 8'hA9,
			8'h00, 8'h38, 8'hE5, 8'h2B, 8'h85, 8'h2B, 8'hA9, 8'h00, 8'hE5, 8'h2C, 8'h85, 8'h2C, 8'h20, 8'h43, 8'hF1, 8'hA9,
			8'h00, 8'h38, 8'hE5, 8'h2E, 8'h85, 8'h2E, 8'hA9, 8'h00, 8'hE5, 8'h2F, 8'h85, 8'h2F, 8'hA9, 8'h00, 8'hE5, 8'h30,
			8'h85, 8'h30, 8'h60, 8'h8A, 8'h48, 8'hA9, 8'h00, 8'h85, 8'h2E, 8'h85, 8'h2F, 8'h85, 8'h30, 8'hA2, 8'h08, 8'h06,
			8'h2E, 8'h26, 8'h2F, 8'h26, 8'h30, 8'h06, 8'h2D, 8'h90, 8'h13, 8'h18, 8'hA5, 8'h2B, 8'h65, 8'h2E, 8'h85, 8'h2E,
			8'hA5, 8'h2C, 8'h65, 8'h2F, 8'h85, 8'h2F, 8'hA9, 8'h00, 8'h65, 8'h30, 8'h85, 8'h30, 8'hCA, 8'hD0, 8'hE0, 8'h68,
			8'hAA, 8'h60, 8'hBD, 8'h24, 8'h04, 8'h85, 8'h2B, 8'hBD, 8'h2D, 8'h04, 8'h85, 8'h2C, 8'hA9, 8'hCD, 8'h20, 8'h19,
			8'hF1, 8'hA5, 8'h2F, 8'h9D, 8'h24, 8'h04, 8'hA5, 8'h30, 8'h9D, 8'h2D, 8'h04, 8'h60, 8'hBD, 8'h12, 8'h04, 8'h85,
			8'h2B, 8'hBD, 8'h1B, 8'h04, 8'h85, 8'h2C, 8'hA9, 8'hCD, 8'h20, 8'h19, 8'hF1, 8'hA5, 8'h2F, 8'h9D, 8'h12, 8'h04,
			8'hA5, 8'h30, 8'h9D, 8'h1B, 8'h04, 8'h60, 8'hA0, 8'h04, 8'hA5, 8'h13, 8'h0A, 8'h66, 8'h13, 8'h66, 8'h12, 8'h88,
			8'hD0, 8'hF6, 8'h60, 8'h8A, 8'h48, 8'hA2, 8'h0B, 8'h06, 8'h1B, 8'h26, 8'h1C, 8'h2A, 8'h2A, 8'h45, 8'h1B, 8'h2A,
			8'h45, 8'h1B, 8'h4A, 8'h4A, 8'h49, 8'hFF, 8'h29, 8'h01, 8'h05, 8'h1B, 8'h85, 8'h1B, 8'hCA, 8'hD0, 8'hE8, 8'h68,
			8'hAA, 8'hA5, 8'h1B, 8'h60, 8'h20, 8'hC1, 8'hDA, 8'hA2, 8'h09, 8'hA9, 8'h00, 8'h95, 8'h03, 8'hCA, 8'h10, 8'hF9,
			8'h85, 8'h3E, 8'hE6, 8'h41, 8'h20, 8'hDE, 8'hD6, 8'hA9, 8'h0F, 8'h8D, 8'h15, 8'h40, 8'hA9, 8'h01, 8'h85, 8'hF0,
			8'hA9, 8'h02, 8'h85, 8'h41, 8'hA4, 8'h40, 8'hD0, 8'h02, 8'hA9, 8'hFF, 8'h85, 8'h42, 8'hA2, 8'h00, 8'h8E, 8'h88,
			8'h04, 8'h86, 8'h3B, 8'h86, 8'h3C, 8'h8E, 8'h58, 8'h05, 8'hCA, 8'h86, 8'h89, 8'hA6, 8'h40, 8'h20, 8'hB0, 8'hF3,
			8'hCA, 8'h10, 8'hFA, 8'hA9, 8'h00, 8'h85, 8'hC8, 8'hA5, 8'h3C, 8'h4A, 8'h4A, 8'hC9, 8'h08, 8'h90, 8'h02, 8'hA9,
			8'h08, 8'hAA, 8'hBD, 8'hBA, 8'hF3, 8'h85, 8'hC6, 8'hBD, 8'hC3, 8'hF3, 8'h85, 8'hC7, 8'hA5, 8'h3C, 8'hC9, 8'h02,
			8'hB0, 8'h06, 8'hA9, 8'h03, 8'h85, 8'hC6, 8'h85, 8'hC7, 8'hA2, 8'h07, 8'hA9, 8'h00, 8'h9D, 8'h48, 8'h04, 8'h9D,
			8'h75, 8'h04, 8'h9D, 8'h7E, 8'h04, 8'h9D, 8'h24, 8'h04, 8'h9D, 8'h2D, 8'h04, 8'h9D, 8'h12, 8'h04, 8'h9D, 8'h1B,
			8'h04, 8'h9D, 8'h63, 8'h04, 8'h9D, 8'h6C, 8'h04, 8'h9D, 8'h00, 8'h04, 8'h9D, 8'h09, 8'h04, 8'hA9, 8'h01, 8'h9D,
			8'h3F, 8'h04, 8'h9D, 8'h5A, 8'h04, 8'hA9, 8'h03, 8'h9D, 8'h36, 8'h04, 8'hCA, 8'h10, 8'hCD, 8'hA2, 8'h05, 8'hA9,
			8'hFF, 8'h95, 8'h8A, 8'hCA, 8'h10, 8'hF9, 8'hA6, 8'h40, 8'h20, 8'h86, 8'hF3, 8'hCA, 8'h10, 8'hFA, 8'h20, 8'h46,
			8'hD2, 8'h20, 8'h93, 8'hD2, 8'hA5, 8'hC6, 8'hC9, 8'h10, 8'hB0, 8'h04, 8'hA9, 8'h58, 8'h85, 8'hC6, 8'h20, 8'hA5,
			8'hF4, 8'h20, 8'hFF, 8'hD8, 8'hA5, 8'h16, 8'hF0, 8'h03, 8'h4C, 8'hC5, 8'hC1, 8'hA5, 8'hC8, 8'hF0, 8'h03, 8'h4C,
			8'h13, 8'hCF, 8'h20, 8'h16, 8'hC7, 8'hA5, 8'h3B, 8'h29, 8'h03, 8'hD0, 8'h08, 8'hA9, 8'h08, 8'h85, 8'hF2, 8'hA6,
			8'h3A, 8'hD0, 8'h06, 8'hA9, 8'hFF, 8'h85, 8'h3D, 8'hE6, 8'h3C, 8'h20, 8'h70, 8'hF4, 8'hA5, 8'h3D, 8'hF0, 8'h05,
			8'hC6, 8'h3D, 8'h20, 8'hCC, 8'hF3, 8'h20, 8'hB3, 8'hF1, 8'h20, 8'h91, 8'hE6, 8'h20, 8'hF9, 8'hC6, 8'h20, 8'h90,
			8'hC7, 8'h20, 8'h31, 8'hC8, 8'h20, 8'hB7, 8'hC8, 8'h20, 8'hDD, 8'hD8, 8'h20, 8'h87, 8'hE5, 8'h20, 8'h74, 8'hCB,
			8'hE6, 8'h4C, 8'hA6, 8'h40, 8'hB5, 8'h88, 8'h10, 8'h25, 8'hA5, 8'h3A, 8'hD0, 8'h3A, 8'hB5, 8'h41, 8'h30, 8'h1D,
			8'hD6, 8'hC3, 8'hD0, 8'h33, 8'h8A, 8'h48, 8'h20, 8'h26, 8'hC7, 8'h68, 8'hAA, 8'hA0, 8'h02, 8'hD6, 8'h41, 8'h84,
			8'h46, 8'h30, 8'h0A, 8'h20, 8'h86, 8'hF3, 8'h20, 8'hB0, 8'hF3, 8'hA9, 8'h80, 8'h85, 8'hF2, 8'hCA, 8'h10, 8'hD4,
			8'hA5, 8'h41, 8'h10, 8'h04, 8'hA5, 8'h42, 8'h30, 8'h4E, 8'hA5, 8'h3A, 8'hF0, 8'h0B, 8'h20, 8'h68, 8'hE7, 8'hAD,
			8'h1C, 8'h06, 8'h29, 8'h30, 8'hF0, 8'h93, 8'h60, 8'hA2, 8'h05, 8'hB5, 8'h8A, 8'hF0, 8'h02, 8'h10, 8'h8A, 8'hCA,
			8'h10, 8'hF7, 8'hA5, 8'hBB, 8'h10, 8'h83, 8'hA6, 8'h40, 8'hB4, 8'h88, 8'h88, 8'h10, 8'h0F, 8'hB5, 8'h41, 8'h30,
			8'h0B, 8'hA9, 8'hFF, 8'h95, 8'h88, 8'hA9, 8'h01, 8'h95, 8'hC3, 8'h4C, 8'hB9, 8'hF2, 8'hCA, 8'h10, 8'hE9, 8'hA9,
			8'h02, 8'h85, 8'hF2, 8'hA2, 8'h96, 8'h20, 8'h5E, 8'hF4, 8'hA6, 8'h3B, 8'hE8, 8'hE0, 8'h10, 8'hD0, 8'h02, 8'hA2,
			8'h04, 8'h86, 8'h3B, 8'h4C, 8'h13, 8'hF2, 8'hA9, 8'h01, 8'h85, 8'hF2, 8'hA9, 8'h00, 8'h85, 8'h17, 8'h85, 8'h18,
			8'h85, 8'h15, 8'h20, 8'h0B, 8'hF4, 8'h20, 8'h65, 8'hF4, 8'h20, 8'h68, 8'hE7, 8'h29, 8'h30, 8'hD0, 8'h04, 8'hC6,
			8'h15, 8'hD0, 8'hF2, 8'h4C, 8'hD4, 8'hF1, 8'hB5, 8'h41, 8'h30, 8'h23, 8'hBD, 8'hAE, 8'hF3, 8'h95, 8'h91, 8'hA9,
			8'hB8, 8'h95, 8'h9A, 8'h95, 8'hBD, 8'hA9, 8'hC8, 8'h95, 8'hBF, 8'hA9, 8'h5A, 8'hB4, 8'h41, 8'h10, 8'h02, 8'hA9,
			8'h01, 8'h95, 8'hC3, 8'hA9, 8'h00, 8'h95, 8'hC1, 8'h9D, 8'h2D, 8'h04, 8'h9D, 8'h24, 8'h04, 8'h60, 8'h20, 8'hD0,
			8'hA9, 8'h03, 8'h9D, 8'h51, 8'h04, 8'hA9, 8'h02, 8'h95, 8'h88, 8'h60, 8'h58, 8'h50, 8'h58, 8'h50, 8'h50, 8'h40,
			8'h38, 8'h30, 8'h28, 8'h04, 8'h04, 8'h03, 8'h03, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'hA5, 8'h3D, 8'h29, 8'h20,
			8'hF0, 8'h1C, 8'hA2, 8'h0A, 8'hBD, 8'hF5, 8'hF3, 8'h95, 8'h57, 8'hCA, 8'h10, 8'hF8, 8'hA0, 8'h0A, 8'hA5, 8'h3C,
			8'h85, 8'h43, 8'h20, 8'h7C, 8'hD7, 8'h85, 8'h60, 8'hA5, 8'h43, 8'h85, 8'h61, 8'h4C, 8'h2D, 8'hC1, 8'hA9, 8'h00,
			8'hA0, 8'hF4, 8'h4C, 8'h31, 8'hC1, 8'h20, 8'h6C, 8'h08, 8'h19, 8'h11, 8'h0A, 8'h1C, 8'h0E, 8'h25, 8'h00, 8'h00,
			8'h20, 8'h6C, 8'h08, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h20, 8'h65, 8'hF4, 8'hA2, 8'h01,
			8'hBD, 8'h3B, 8'hF4, 8'hBC, 8'h3D, 8'hF4, 8'h20, 8'h31, 8'hC1, 8'hCA, 8'h10, 8'hF4, 8'hA2, 8'h0F, 8'hA9, 8'h24,
			8'h95, 8'h5A, 8'hCA, 8'h10, 8'hF9, 8'hA9, 8'h10, 8'h85, 8'h59, 8'hA9, 8'h21, 8'h85, 8'h57, 8'hA2, 8'h02, 8'hBD,
			8'h3F, 8'hF4, 8'h85, 8'h58, 8'h20, 8'h2D, 8'hC1, 8'hCA, 8'h10, 8'hF5, 8'h60, 8'h42, 8'h55, 8'hF4, 8'hF4, 8'h88,
			8'hA8, 8'hE8, 8'h21, 8'hC8, 8'h10, 8'h24, 8'h24, 8'h24, 8'h10, 8'h0A, 8'h16, 8'h0E, 8'h24, 8'h24, 8'h18, 8'h1F,
			8'h0E, 8'h1B, 8'h24, 8'h24, 8'h24, 8'h23, 8'hDA, 8'h04, 8'hAA, 8'hAA, 8'hAA, 8'hAA, 8'hA2, 8'h14, 8'h20, 8'h65,
			8'hF4, 8'hCA, 8'hD0, 8'hFA, 8'h60, 8'hA9, 8'h00, 8'h85, 8'h02, 8'hA5, 8'h02, 8'hF0, 8'hFC, 8'hC6, 8'h02, 8'h60,
			8'h20, 8'h69, 8'hF4, 8'hA5, 8'h3A, 8'hD0, 8'hF8, 8'h20, 8'h68, 8'hE7, 8'h29, 8'h10, 8'hF0, 8'hF1, 8'hA9, 8'h04,
			8'h85, 8'hF2, 8'hA5, 8'h01, 8'h29, 8'hEF, 8'h8D, 8'h01, 8'h20, 8'h20, 8'h65, 8'hF4, 8'h20, 8'h68, 8'hE7, 8'h29,
			8'h10, 8'hF0, 8'hF6, 8'hA5, 8'h01, 8'h8D, 8'h01, 8'h20, 8'hA0, 8'h04, 8'hA5, 8'hC8, 8'h05, 8'h16, 8'hF0, 8'h02,
			8'hA0, 8'h20, 8'h84, 8'hF2, 8'h60, 8'hA9, 8'h01, 8'h8D, 8'h8E, 8'h04, 8'h8D, 8'h8F, 8'h04, 8'hA9, 8'hFF, 8'h85,
			8'hBB, 8'h85, 8'h87, 8'h8D, 8'h8C, 8'h04, 8'hA2, 8'h01, 8'h8E, 8'h59, 8'h04, 8'h86, 8'h90, 8'hE8, 8'h86, 8'h46,
			8'hA9, 8'h40, 8'h85, 8'h99, 8'h60, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'h20, 8'h8F, 8'hF7, 8'h60, 8'hA9, 8'h00, 8'hAA, 8'h85, 8'hFD, 8'hF0, 8'h10, 8'h8A, 8'h4A, 8'hAA, 8'hE8, 8'h8A,
			8'hC9, 8'h04, 8'hF0, 8'hEF, 8'hA5, 8'hFD, 8'h18, 8'h69, 8'h04, 8'h85, 8'hFD, 8'h8A, 8'h0A, 8'hAA, 8'hB5, 8'hE0,
			8'h85, 8'hFE, 8'hB5, 8'hE1, 8'h85, 8'hFF, 8'hB5, 8'hE1, 8'hF0, 8'hE1, 8'h8A, 8'h4A, 8'hAA, 8'hD6, 8'hD0, 8'hD0,
			8'hDD, 8'hB4, 8'hE8, 8'hF6, 8'hE8, 8'hB1, 8'hFE, 8'hF0, 8'hC7, 8'hA8, 8'hC9, 8'hFF, 8'hF0, 8'h09, 8'h29, 8'hC0,
			8'hC9, 8'hC0, 8'hF0, 8'h0F, 8'h4C, 8'h61, 8'hF5, 8'hB5, 8'hD8, 8'hF0, 8'h13, 8'hD6, 8'hD8, 8'hB5, 8'hEC, 8'h95,
			8'hE8, 8'hD0, 8'h0B, 8'h98, 8'h29, 8'h3F, 8'h95, 8'hD8, 8'hD6, 8'hD8, 8'hB5, 8'hE8, 8'h95, 8'hEC, 8'h4C, 8'h31,
			8'hF5, 8'h98, 8'h10, 8'h17, 8'h29, 8'h0F, 8'h18, 8'h65, 8'hDF, 8'hA8, 8'hB9, 8'h60, 8'hF6, 8'h95, 8'hD4, 8'hA8,
			8'h8A, 8'hC9, 8'h02, 8'hF0, 8'h4F, 8'hB4, 8'hE8, 8'hF6, 8'hE8, 8'hB1, 8'hFE, 8'hA8, 8'h8A, 8'hC9, 8'h03, 8'hF0,
			8'h60, 8'h48, 8'hAA, 8'hC9, 8'h01, 8'hF0, 8'h32, 8'hA6, 8'hFD, 8'hB9, 8'h01, 8'hF6, 8'hF0, 8'h0B, 8'h9D, 8'h02,
			8'h40, 8'hB9, 8'h00, 8'hF6, 8'h09, 8'h08, 8'h9D, 8'h03, 8'h40, 8'hA8, 8'h68, 8'hAA, 8'h98, 8'hD0, 8'h0B, 8'hA0,
			8'h00, 8'h8A, 8'hC9, 8'h02, 8'hF0, 8'h06, 8'hA0, 8'h10, 8'hD0, 8'h02, 8'hB4, 8'hDC, 8'h98, 8'hA4, 8'hFD, 8'h99,
			8'h00, 8'h40, 8'hB5, 8'hD4, 8'h95, 8'hD0, 8'h4C, 8'h0E, 8'hF5, 8'hA5, 8'hF5, 8'h29, 8'h02, 8'hF0, 8'hC8, 8'h68,
			8'hAA, 8'h4C, 8'hB2, 8'hF5, 8'h98, 8'hAC, 8'hF0, 8'h07, 8'hF0, 8'h04, 8'hA9, 8'hFF, 8'hD0, 8'h0B, 8'h18, 8'h69,
			8'hFE, 8'h0A, 8'h0A, 8'hC9, 8'h3C, 8'h90, 8'h02, 8'hA9, 8'h3C, 8'h8D, 8'h08, 8'h40, 8'h85, 8'hDE, 8'h4C, 8'h75,
			8'hF5, 8'hA5, 8'hF4, 8'hC9, 8'h02, 8'hF0, 8'h12, 8'hB9, 8'h00, 8'hF7, 8'h8D, 8'h0C, 8'h40, 8'hB9, 8'h01, 8'hF7,
			8'h8D, 8'h0E, 8'h40, 8'hB9, 8'h02, 8'hF7, 8'h8D, 8'h0F, 8'h40, 8'h4C, 8'hB2, 8'hF5, 8'h16, 8'hFF, 8'h10, 8'hC5,
			8'h07, 8'hF0, 8'h00, 8'h00, 8'h00, 8'hD4, 8'h00, 8'hC8, 8'h00, 8'hBD, 8'h00, 8'hB2, 8'h00, 8'hA8, 8'h00, 8'h9F,
			8'h00, 8'h96, 8'h00, 8'h8D, 8'h00, 8'h85, 8'h00, 8'h7E, 8'h00, 8'h76, 8'h00, 8'h70, 8'h01, 8'hAB, 8'h01, 8'h93,
			8'h01, 8'h7C, 8'h01, 8'h67, 8'h01, 8'h52, 8'h01, 8'h3F, 8'h01, 8'h2D, 8'h01, 8'h1C, 8'h01, 8'h0C, 8'h00, 8'hFD,
			8'h00, 8'hEE, 8'h00, 8'hE1, 8'h03, 8'h57, 8'h03, 8'h27, 8'h02, 8'hF9, 8'h02, 8'hCF, 8'h02, 8'hA6, 8'h02, 8'h80,
			8'h02, 8'h5C, 8'h02, 8'h3A, 8'h02, 8'h1A, 8'h01, 8'hFC, 8'h01, 8'hDF, 8'h01, 8'hC4, 8'h03, 8'hF8, 8'h00, 8'h69,
			8'h00, 8'h63, 8'h00, 8'h5E, 8'h00, 8'h58, 8'h00, 8'h53, 8'h00, 8'h4F, 8'h00, 8'h4A, 8'h00, 8'h46, 8'h00, 8'h42,
			8'h03, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h12, 8'h24, 8'h09, 8'h08, 8'h04, 8'h07, 8'h01, 8'h04, 8'h08, 8'h10, 8'h20,
			8'h40, 8'h18, 8'h30, 8'h0C, 8'h01, 8'h06, 8'h0C, 8'h18, 8'h30, 8'h60, 8'h24, 8'h48, 8'h12, 8'h10, 8'h08, 8'h0E,
			8'h02, 8'h03, 8'h04, 8'hA9, 8'h00, 8'hF0, 8'h0A, 8'hA9, 8'h08, 8'hD0, 8'h06, 8'hA9, 8'h0C, 8'hD0, 8'h02, 8'hA9,
			8'h04, 8'h85, 8'hF9, 8'hA9, 8'h40, 8'h85, 8'hFA, 8'h86, 8'hFB, 8'h84, 8'hFC, 8'hA0, 8'h00, 8'hB1, 8'hFB, 8'h91,
			8'hF9, 8'hC8, 8'h98, 8'hC9, 8'h04, 8'hD0, 8'hF6, 8'h60, 8'hAA, 8'h20, 8'h98, 8'hF7, 8'h86, 8'hF6, 8'hAD, 8'hF5,
			8'h07, 8'hF0, 8'h0B, 8'hC9, 8'h02, 8'hD0, 8'h07, 8'h85, 8'hF0, 8'hA9, 8'h00, 8'h8D, 8'hF5, 8'h07, 8'hB9, 8'hCA,
			8'hFB, 8'hA8, 8'hA2, 8'h00, 8'hB9, 8'hCA, 8'hFB, 8'h95, 8'hDF, 8'hC8, 8'hE8, 8'h8A, 8'hC9, 8'h09, 8'hD0, 8'hF4,
			8'hA9, 8'h01, 8'h85, 8'hD0, 8'h85, 8'hD1, 8'h85, 8'hD2, 8'h85, 8'hD3, 8'hA9, 8'h00, 8'h85, 8'hE8, 8'h85, 8'hE9,
			8'h85, 8'hEA, 8'h85, 8'hEB, 8'h60, 8'h94, 8'hAB, 8'hFD, 8'h58, 8'h00, 8'h7F, 8'h04, 8'h18, 8'h3F, 8'h7F, 8'h00,
			8'h00, 8'h06, 8'h7F, 8'h0A, 8'hC0, 8'h08, 8'h7F, 8'h05, 8'hC0, 8'hC1, 8'h89, 8'h02, 8'h0F, 8'hFF, 8'hFF, 8'hFF,
			8'h10, 8'h00, 8'h18, 8'h10, 8'h01, 8'h18, 8'h00, 8'h01, 8'h88, 8'h02, 8'h02, 8'h40, 8'h03, 8'h05, 8'h40, 8'h04,
			8'h07, 8'h40, 8'hA9, 8'h7F, 8'h8D, 8'h01, 8'h40, 8'h8D, 8'h05, 8'h40, 8'h86, 8'hDC, 8'h84, 8'hDD, 8'h60, 8'hA2,
			8'hE5, 8'hA0, 8'hF6, 8'hD0, 8'h20, 8'hA5, 8'hF3, 8'h4A, 8'hB0, 8'h0C, 8'hA5, 8'hF7, 8'h4A, 8'hB0, 8'h1A, 8'hA5,
			8'hF0, 8'h29, 8'h10, 8'hD0, 8'hEA, 8'h60, 8'hA5, 8'hF7, 8'h09, 8'h01, 8'h85, 8'hF7, 8'hA9, 8'h00, 8'h8D, 8'hE4,
			8'h07, 8'hA2, 8'hFC, 8'hA0, 8'hF5, 8'h20, 8'h83, 8'hF6, 8'h60, 8'hEE, 8'hE4, 8'h07, 8'hAD, 8'hE4, 8'h07, 8'hC9,
			8'h58, 8'hD0, 8'h28, 8'hA9, 8'h00, 8'h85, 8'hF7, 8'h60, 8'hA9, 8'hC0, 8'h8D, 8'h17, 8'h40, 8'h20, 8'h25, 8'hFB,
			8'h20, 8'h0A, 8'hF9, 8'h20, 8'h38, 8'hFA, 8'h20, 8'hAC, 8'hFA, 8'h20, 8'h24, 8'hF8, 8'hA5, 8'hF1, 8'h8D, 8'hE9,
			8'h07, 8'hA9, 8'h00, 8'h85, 8'hF0, 8'h85, 8'hF1, 8'h85, 8'hF2, 8'h85, 8'hF3, 8'h60, 8'hA5, 8'hF4, 8'h29, 8'h06,
			8'hD0, 8'hF9, 8'hA5, 8'hF4, 8'h29, 8'hF0, 8'h85, 8'hF4, 8'hA2, 8'hE9, 8'hA0, 8'hF6, 8'h4C, 8'h79, 8'hF8, 8'hA5,
			8'hF6, 8'hC9, 8'h20, 8'hD0, 8'h0A, 8'hEE, 8'hE8, 8'h07, 8'h29, 8'h0F, 8'hC9, 8'h0F, 8'hD0, 8'h07, 8'h8A, 8'hA5,
			8'hF4, 8'h29, 8'h20, 8'hD0, 8'h22, 8'hA9, 8'h10, 8'h8D, 8'h0C, 8'h40, 8'h8D, 8'h00, 8'h40, 8'h8D, 8'h04, 8'h40,
			8'hA9, 8'h00, 8'h85, 8'hF4, 8'h85, 8'hF5, 8'h85, 8'hF6, 8'h8D, 8'hFA, 8'h07, 8'h85, 8'hF7, 8'h8D, 8'h08, 8'h40,
			8'h8D, 8'h11, 8'h40, 8'h8D, 8'hF0, 8'h07, 8'h60, 8'hA9, 8'h10, 8'h8D, 8'h04, 8'h40, 8'h8D, 8'h0C, 8'h40, 8'hA9,
			8'h00, 8'hF0, 8'hE1, 8'hA9, 8'h00, 8'h8D, 8'hFA, 8'h07, 8'h60, 8'hA2, 8'hF5, 8'hA0, 8'hF6, 8'h4C, 8'h79, 8'hF8,
			8'hEE, 8'hFB, 8'h07, 8'hAD, 8'hFB, 8'h07, 8'hC9, 8'h10, 8'hF0, 8'hEF, 8'hC9, 8'h20, 8'hF0, 8'hE5, 8'h60, 8'hA9,
			8'h00, 8'h8D, 8'hFB, 8'h07, 8'hA9, 8'hF0, 8'h8D, 8'hFA, 8'h07, 8'hA2, 8'hF1, 8'hA0, 8'hF6, 8'h4C, 8'h79, 8'hF8,
			8'hA5, 8'hF4, 8'h29, 8'hF0, 8'h09, 8'h02, 8'h85, 8'hF4, 8'hA9, 8'h00, 8'h8D, 8'hF7, 8'h07, 8'hA2, 8'hF1, 8'hA0,
			8'hF6, 8'h4C, 8'h79, 8'hF8, 8'hEE, 8'hF7, 8'h07, 8'hAD, 8'hF7, 8'h07, 8'hC9, 8'h10, 8'hD0, 8'h3D, 8'h4C, 8'h9B,
			8'hF8, 8'h4C, 8'hA5, 8'hF7, 8'hA5, 8'hF0, 8'h4A, 8'hB0, 8'hF8, 8'hA5, 8'hF6, 8'hC9, 8'hDF, 8'hF0, 8'h0C, 8'hC9,
			8'h7F, 8'hF0, 8'h08, 8'hC9, 8'h20, 8'hF0, 8'h04, 8'hA5, 8'hF6, 8'hD0, 8'h20, 8'hAD, 8'hFA, 8'h07, 8'hC9, 8'h0F,
			8'hF0, 8'hAD, 8'hC9, 8'hF0, 8'hF0, 8'h9A, 8'hA5, 8'hF0, 8'h4A, 8'h4A, 8'hB0, 8'hB4, 8'h4A, 8'hB0, 8'h10, 8'h4A,
			8'hB0, 8'h0A, 8'hA5, 8'hF4, 8'h4A, 8'h4A, 8'hB0, 8'hBC, 8'h4A, 8'hB0, 8'h22, 8'h60, 8'h4C, 8'h7C, 8'hF7, 8'hA5,
			8'hF4, 8'h29, 8'h80, 8'hD0, 8'hF6, 8'hA5, 8'hF4, 8'h29, 8'hF0, 8'h09, 8'h04, 8'h85, 8'hF4, 8'hA9, 8'h00, 8'h8D,
			8'hF3, 8'h07, 8'h8D, 8'hF1, 8'h07, 8'hA2, 8'hED, 8'hA0, 8'hF6, 8'h20, 8'h8B, 8'hF6, 8'h60, 8'hEE, 8'hF3, 8'h07,
			8'hAD, 8'hF3, 8'h07, 8'hC9, 8'h03, 8'hD0, 8'h1A, 8'hA9, 8'h00, 8'h8D, 8'hF3, 8'h07, 8'hEE, 8'hF1, 8'h07, 8'hAD,
			8'hF1, 8'h07, 8'hC9, 8'h10, 8'hD0, 8'h0C, 8'hA9, 8'h10, 8'h8D, 8'h0C, 8'h40, 8'hA5, 8'hF4, 8'h29, 8'hF0, 8'h85,
			8'hF4, 8'h60, 8'h8D, 8'h0E, 8'h40, 8'h60, 8'hA9, 8'h00, 8'h8D, 8'hE0, 8'h07, 8'h18, 8'hA5, 8'h1B, 8'h29, 8'h07,
			8'h69, 8'h02, 8'h8D, 8'hE1, 8'h07, 8'hA5, 8'hF7, 8'h29, 8'h00, 8'h09, 8'h80, 8'h85, 8'hF7, 8'hD0, 8'h29, 8'hEE,
			8'hE0, 8'h07, 8'hAD, 8'hE0, 8'h07, 8'hCD, 8'hE1, 8'h07, 8'hD0, 8'h1E, 8'hA9, 8'h10, 8'h8D, 8'h00, 8'h40, 8'h8D,
			8'h04, 8'h40, 8'hA9, 8'h00, 8'h85, 8'hF7, 8'hA5, 8'hF4, 8'h29, 8'h0F, 8'h85, 8'hF4, 8'h60, 8'h20, 8'hA5, 8'hF7,
			8'hA9, 8'h80, 8'h85, 8'hF4, 8'hA9, 8'h02, 8'h85, 8'hF0, 8'hA2, 8'hF9, 8'hA0, 8'hF6, 8'h20, 8'h83, 8'hF6, 8'hA5,
			8'h1B, 8'h29, 8'h0F, 8'h8D, 8'h02, 8'h40, 8'hA2, 8'hF9, 8'hA0, 8'hF6, 8'h20, 8'h8F, 8'hF6, 8'hA5, 8'h1B, 8'h4A,
			8'h4A, 8'h29, 8'h0F, 8'h8D, 8'h06, 8'h40, 8'h60, 8'h4C, 8'hA6, 8'hF8, 8'hA5, 8'hF6, 8'hF0, 8'h0D, 8'hC9, 8'hDF,
			8'hF0, 8'h09, 8'hA5, 8'hF0, 8'h29, 8'hE0, 8'hF0, 8'h36, 8'h20, 8'hA5, 8'hF7, 8'hA5, 8'hF0, 8'h0A, 8'hB0, 8'hBD,
			8'h0A, 8'hB0, 8'h2F, 8'h0A, 8'hB0, 8'h3F, 8'hA5, 8'hF4, 8'h0A, 8'hB0, 8'hBD, 8'hA5, 8'hF4, 8'h29, 8'hE0, 8'hD0,
			8'h1D, 8'hA5, 8'hF6, 8'hC9, 8'hDF, 8'hF0, 8'h14, 8'hA5, 8'hF6, 8'hD0, 8'h13, 8'hA5, 8'hF3, 8'h0A, 8'hB0, 8'hC7,
			8'h0A, 8'hB0, 8'h34, 8'hA5, 8'hF7, 8'h0A, 8'hB0, 8'h07, 8'h0A, 8'hB0, 8'h48, 8'h20, 8'h25, 8'hF7, 8'h60, 8'h4C,
			8'hBF, 8'hF8, 8'hA9, 8'h0F, 8'h8D, 8'hFA, 8'h07, 8'hA5, 8'hF4, 8'h29, 8'h0F, 8'h09, 8'h40, 8'h85, 8'hF4, 8'hA2,
			8'hD1, 8'hA0, 8'hF9, 8'hD0, 8'h2A, 8'hA9, 8'h02, 8'h85, 8'hF0, 8'hA5, 8'hF4, 8'h29, 8'h0F, 8'h09, 8'h20, 8'h85,
			8'hF4, 8'hA2, 8'hCD, 8'hA0, 8'hF9, 8'hD0, 8'h18, 8'hA9, 8'h00, 8'h8D, 8'hFC, 8'h07, 8'hA5, 8'hF7, 8'h29, 8'h00,
			8'h09, 8'h40, 8'h85, 8'hF7, 8'hA2, 8'hD5, 8'hA0, 8'hF9, 8'h20, 8'h8F, 8'hF6, 8'hA2, 8'hD9, 8'hA0, 8'hF9, 8'h20,
			8'h83, 8'hF6, 8'h60, 8'hEE, 8'hFC, 8'h07, 8'hAD, 8'hFC, 8'h07, 8'hC9, 8'h12, 8'hF0, 8'h2D, 8'hC9, 8'h06, 8'h90,
			8'h10, 8'hA5, 8'h1B, 8'h09, 8'h10, 8'h29, 8'h7F, 8'h8D, 8'hFE, 8'h07, 8'h2A, 8'h8D, 8'hFD, 8'h07, 8'h4C, 8'hBD,
			8'hF9, 8'hEE, 8'hFD, 8'h07, 8'hEE, 8'hFD, 8'h07, 8'hEE, 8'hFE, 8'h07, 8'hEE, 8'hFE, 8'h07, 8'hAD, 8'hFD, 8'h07,
			8'h8D, 8'h06, 8'h40, 8'hAD, 8'hFE, 8'h07, 8'h8D, 8'h02, 8'h40, 8'h60, 8'h4C, 8'hCA, 8'hF8, 8'hB8, 8'hD5, 8'h20,
			8'h00, 8'h9F, 8'h93, 8'h80, 8'h22, 8'h3F, 8'hBA, 8'hE0, 8'h06, 8'h3F, 8'hBB, 8'hCE, 8'h06, 8'hB8, 8'h93, 8'h50,
			8'h02, 8'h80, 8'h7F, 8'h60, 8'h68, 8'h80, 8'h7F, 8'h62, 8'h68, 8'hA5, 8'hF5, 8'h29, 8'h02, 8'hD0, 8'h37, 8'hA5,
			8'hF6, 8'hC9, 8'hDF, 8'hF0, 8'h04, 8'hA5, 8'hF6, 8'hD0, 8'h2D, 8'hA9, 8'h00, 8'h8D, 8'hF9, 8'h07, 8'hA5, 8'hF5,
			8'h29, 8'hE0, 8'h09, 8'h02, 8'h85, 8'hF5, 8'hA2, 8'hDD, 8'hA0, 8'hF9, 8'hD0, 8'h73, 8'hEE, 8'hF9, 8'h07, 8'hAD,
			8'hF9, 8'h07, 8'hC9, 8'h07, 8'hD0, 8'h10, 8'hA9, 8'h7F, 8'h8D, 8'h05, 8'h40, 8'hA9, 8'h10, 8'h8D, 8'h04, 8'h40,
			8'hA5, 8'hF5, 8'h29, 8'hE0, 8'h85, 8'hF5, 8'h60, 8'h20, 8'hA5, 8'hF7, 8'hA2, 8'hE1, 8'hA0, 8'hF9, 8'h20, 8'h83,
			8'hF6, 8'hA2, 8'hE5, 8'hA0, 8'hF9, 8'h4C, 8'h7F, 8'hFA, 8'hA5, 8'hF6, 8'hF0, 8'h06, 8'h29, 8'h0F, 8'hC9, 8'h0F,
			8'hD0, 8'h21, 8'hA5, 8'hF4, 8'h29, 8'h80, 8'hD0, 8'h1B, 8'hA5, 8'hF7, 8'h29, 8'hC0, 8'hD0, 8'h15, 8'hA5, 8'hF1,
			8'h4A, 8'hB0, 8'hD4, 8'h4A, 8'hB0, 8'h93, 8'h4A, 8'hB0, 8'h2A, 8'h4A, 8'h4A, 8'hB0, 8'h07, 8'hA5, 8'hF5, 8'h4A,
			8'h4A, 8'hB0, 8'hA9, 8'h60, 8'hA5, 8'hF6, 8'hD0, 8'hFB, 8'hA5, 8'hF5, 8'h29, 8'h02, 8'hD0, 8'hF5, 8'hA2, 8'h8A,
			8'hA0, 8'hFA, 8'h20, 8'h8F, 8'hF6, 8'hA5, 8'h1B, 8'h29, 8'h3F, 8'h09, 8'h10, 8'h8D, 8'h06, 8'h40, 8'h60, 8'h20,
			8'h8F, 8'hF6, 8'h60, 8'hA0, 8'h0A, 8'hA9, 8'hEF, 8'h4C, 8'hA5, 8'hFB, 8'hD9, 8'h86, 8'hA8, 8'h48, 8'h08, 8'h7F,
			8'h40, 8'h28, 8'h08, 8'h7F, 8'h45, 8'h28, 8'hEE, 8'hF6, 8'h07, 8'hAD, 8'hF6, 8'h07, 8'hC9, 8'h04, 8'hD0, 8'h38,
			8'hA5, 8'hF5, 8'h29, 8'h1F, 8'h85, 8'hF5, 8'hA2, 8'h92, 8'hA0, 8'hFA, 8'hD0, 8'h54, 8'hA5, 8'hF6, 8'hF0, 8'h0A,
			8'hC9, 8'h08, 8'hF0, 8'h06, 8'h29, 8'h0F, 8'hC9, 8'h0F, 8'hD0, 8'h1E, 8'hA5, 8'hF4, 8'h29, 8'h80, 8'hD0, 8'h18,
			8'hA5, 8'hF1, 8'h0A, 8'hB0, 8'h52, 8'h0A, 8'hB0, 8'h1A, 8'hA5, 8'hF5, 8'h0A, 8'h0A, 8'hB0, 8'hC8, 8'hA5, 8'hF1,
			8'h29, 8'h20, 8'hF0, 8'h05, 8'hA5, 8'hF6, 8'hF0, 8'h2C, 8'h60, 8'hA5, 8'hF6, 8'hC9, 8'hDF, 8'hD0, 8'hF9, 8'h4C,
			8'h9F, 8'hF7, 8'hA5, 8'hF5, 8'h29, 8'h1F, 8'h09, 8'h40, 8'h85, 8'hF5, 8'hA9, 8'h00, 8'h8D, 8'h08, 8'h40, 8'h85,
			8'hF6, 8'h8D, 8'hF6, 8'h07, 8'hA9, 8'h10, 8'h8D, 8'h04, 8'h40, 8'h8D, 8'h0C, 8'h40, 8'hA2, 8'h8E, 8'hA0, 8'hFA,
			8'h20, 8'h87, 8'hF6, 8'h60, 8'hAD, 8'hE9, 8'h07, 8'h29, 8'h20, 8'hD0, 8'h05, 8'hA9, 8'h02, 8'h8D, 8'hF5, 8'h07,
			8'hA0, 8'h08, 8'hA9, 8'hDF, 8'h4C, 8'hA5, 8'hFB, 8'hA0, 8'h04, 8'hA9, 8'h7F, 8'h4C, 8'hA5, 8'hFB, 8'hA0, 8'h00,
			8'hA9, 8'h02, 8'h4C, 8'hC1, 8'hFB, 8'hAD, 8'hE8, 8'h07, 8'hD0, 8'h34, 8'hA5, 8'hF2, 8'h4A, 8'hB0, 8'h53, 8'h4A,
			8'hB0, 8'hEC, 8'h4A, 8'hB0, 8'h17, 8'h4A, 8'hB0, 8'h44, 8'h4A, 8'hB0, 8'h2E, 8'h4A, 8'hB0, 8'h20, 8'h4A, 8'hB0,
			8'h17, 8'h4A, 8'hB0, 8'h0E, 8'hA5, 8'hF6, 8'hD0, 8'h01, 8'h60, 8'h4C, 8'h04, 8'hF5, 8'hA0, 8'h02, 8'hA9, 8'h04,
			8'hD0, 8'h53, 8'hA0, 8'h09, 8'hA9, 8'h80, 8'hD0, 8'h15, 8'hA0, 8'h07, 8'hA9, 8'h40, 8'hD0, 8'h0F, 8'hA9, 8'h00,
			8'h8D, 8'hE8, 8'h07, 8'hA0, 8'h06, 8'hA9, 8'h20, 8'hD0, 8'h58, 8'hA0, 8'h05, 8'hA9, 8'h10, 8'h20, 8'hA8, 8'hF6,
			8'hA2, 8'hFC, 8'hA0, 8'hFC, 8'h20, 8'h12, 8'hF7, 8'hEE, 8'hF0, 8'h07, 8'hD0, 8'hCD, 8'hA0, 8'h03, 8'hA9, 8'h08,
			8'hD0, 8'h04, 8'hA0, 8'h01, 8'hA9, 8'h01, 8'h20, 8'hA8, 8'hF6, 8'hA2, 8'h80, 8'hA0, 8'h80, 8'h20, 8'h1A, 8'hF7,
			8'hA9, 8'h83, 8'h8D, 8'h01, 8'h40, 8'hA9, 8'h7F, 8'h8D, 8'h05, 8'h40, 8'hD0, 8'h13, 8'h20, 8'hA8, 8'hF6, 8'hA2,
			8'h04, 8'hA0, 8'h04, 8'hD0, 8'h07, 8'h20, 8'hA8, 8'hF6, 8'hA2, 8'h80, 8'hA0, 8'h80, 8'h20, 8'h12, 8'hF7, 8'hA9,
			8'h00, 8'h8D, 8'hF0, 8'h07, 8'hA5, 8'hF4, 8'h29, 8'h20, 8'hF0, 8'h8F, 8'hA9, 8'hD5, 8'h8D, 8'h01, 8'h40, 8'hD0,
			8'h88, 8'h20, 8'hA8, 8'hF6, 8'hA2, 8'h80, 8'hA0, 8'hBA, 8'hD0, 8'hC3, 8'h0B, 8'h14, 8'h1D, 8'h26, 8'h2F, 8'h38,
			8'h41, 8'h4A, 8'h53, 8'h5C, 8'h65, 8'h0C, 8'h02, 8'hFF, 8'h0B, 8'hFF, 8'h1E, 8'hFF, 8'h31, 8'hFF, 8'h15, 8'h18,
			8'hFE, 8'h2A, 8'hFE, 8'h65, 8'hFE, 8'h86, 8'hFE, 8'h0C, 8'h0D, 8'hFE, 8'h00, 8'h00, 8'h13, 8'hFE, 8'h00, 8'h00,
			8'h15, 8'h38, 8'hFF, 8'h5A, 8'hFF, 8'h79, 8'hFF, 8'h94, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hD7, 8'hFE, 8'hED, 8'hFE,
			8'h00, 8'h00, 8'h00, 8'hB3, 8'hFF, 8'hC9, 8'hFF, 8'hDA, 8'hFF, 8'hEF, 8'hFF, 8'h15, 8'hA5, 8'hFC, 8'h0A, 8'hFD,
			8'h98, 8'hFD, 8'hE0, 8'hFD, 8'h15, 8'hB2, 8'hFE, 8'h00, 8'h00, 8'hC5, 8'hFE, 8'h00, 8'h00, 8'h15, 8'h00, 8'h00,
			8'h92, 8'hFE, 8'hA1, 8'hFE, 8'h00, 8'h00, 8'h0C, 8'h59, 8'hFC, 8'h72, 8'hFC, 8'h8C, 8'hFC, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h38, 8'hFC, 8'h49, 8'hFC, 8'h00, 8'h00, 8'h82, 8'h02, 8'h8B, 8'h02, 8'h80, 8'h08, 8'h02, 8'h10,
			8'h02, 8'h16, 8'h02, 8'h52, 8'h02, 8'h02, 8'h02, 8'h1A, 8'h00, 8'h82, 8'h02, 8'h80, 8'h10, 8'h02, 8'h16, 8'h02,
			8'h52, 8'h02, 8'h5A, 8'h02, 8'h02, 8'h02, 8'h56, 8'h81, 8'h02, 8'h80, 8'h12, 8'h02, 8'h0C, 8'h02, 8'h04, 8'h02,
			8'h0C, 8'h02, 8'h04, 8'h02, 8'h2A, 8'h02, 8'h81, 8'h04, 8'h02, 8'h80, 8'h04, 8'h02, 8'h81, 8'h04, 8'h88, 8'h02,
			8'h02, 8'h00, 8'h88, 8'h02, 8'h02, 8'h80, 8'h04, 8'h02, 8'h2A, 8'h02, 8'h24, 8'h02, 8'h2A, 8'h02, 8'h24, 8'h02,
			8'h1C, 8'h02, 8'h81, 8'h22, 8'h02, 8'h80, 8'h22, 8'h02, 8'h81, 8'h24, 8'h88, 8'h02, 8'h88, 8'h02, 8'h80, 8'h56,
			8'h02, 8'h4E, 8'h02, 8'h12, 8'h02, 8'h4E, 8'h02, 8'h12, 8'h02, 8'h0C, 8'h02, 8'h81, 8'h10, 8'h02, 8'h80, 8'h10,
			8'h02, 8'h81, 8'h12, 8'h88, 8'h02, 8'hC3, 8'h81, 8'h02, 8'h02, 8'h1C, 8'h02, 8'h02, 8'h02, 8'h1C, 8'h1C, 8'hFF,
			8'hC6, 8'h88, 8'h1C, 8'hFF, 8'hC7, 8'h82, 8'h4C, 8'h4C, 8'h2A, 8'h4C, 8'hFF, 8'hC6, 8'h88, 8'h1C, 8'hFF, 8'hC4,
			8'h81, 8'h46, 8'h02, 8'h46, 8'h02, 8'h32, 8'h02, 8'h46, 8'h80, 8'h2E, 8'h2E, 8'hFF, 8'hC3, 8'h82, 8'h46, 8'h46,
			8'h81, 8'h32, 8'h32, 8'h46, 8'h2E, 8'hFF, 8'h80, 8'h0C, 8'h0C, 8'h81, 8'h46, 8'h46, 8'h46, 8'h80, 8'h04, 8'h04,
			8'h81, 8'h46, 8'h46, 8'h02, 8'hC8, 8'h82, 8'h4C, 8'h4C, 8'h2A, 8'h4C, 8'hFF, 8'hC2, 8'h81, 8'h46, 8'h80, 8'h32,
			8'h32, 8'h82, 8'h46, 8'h04, 8'h81, 8'h46, 8'h2A, 8'hFF, 8'hC2, 8'h81, 8'h0C, 8'h0C, 8'h80, 8'h04, 8'h04, 8'h81,
			8'h04, 8'h80, 8'h2E, 8'h2E, 8'h81, 8'h2E, 8'h82, 8'h24, 8'hFF, 8'h00, 8'h81, 8'h32, 8'h02, 8'h02, 8'h06, 8'h0C,
			8'h32, 8'h02, 8'h02, 8'h8A, 8'h2E, 8'h8B, 8'h02, 8'h8A, 8'h2E, 8'h8B, 8'h02, 8'h8A, 8'h2E, 8'h8B, 8'h02, 8'h88,
			8'h2E, 8'h32, 8'h2E, 8'hD0, 8'h8C, 8'h2C, 8'h24, 8'hFF, 8'hD0, 8'h2E, 8'h20, 8'hFF, 8'hC3, 8'h80, 8'h28, 8'h02,
			8'h82, 8'h02, 8'h80, 8'h2C, 8'h02, 8'h32, 8'h02, 8'h24, 8'h02, 8'h82, 8'h02, 8'h81, 8'h02, 8'h80, 8'h28, 8'h02,
			8'h06, 8'h02, 8'h28, 8'h02, 8'h81, 8'h02, 8'h80, 8'h24, 8'h02, 8'h32, 8'h02, 8'h24, 8'h02, 8'hFF, 8'h80, 8'h28,
			8'h02, 8'h82, 8'h02, 8'h80, 8'h2C, 8'h02, 8'h32, 8'h02, 8'h24, 8'h02, 8'h82, 8'h02, 8'h89, 8'h0C, 8'h0A, 8'h08,
			8'h06, 8'h32, 8'h30, 8'h2E, 8'h2C, 8'h2A, 8'h28, 8'h26, 8'h24, 8'h02, 8'h02, 8'h02, 8'h86, 8'h02, 8'hC7, 8'h84,
			8'h02, 8'hFF, 8'hC4, 8'h80, 8'h28, 8'h02, 8'h82, 8'h02, 8'h80, 8'h2C, 8'h02, 8'h32, 8'h02, 8'h24, 8'h02, 8'h82,
			8'h02, 8'h81, 8'h02, 8'h80, 8'h28, 8'h02, 8'h06, 8'h02, 8'h28, 8'h02, 8'h81, 8'h02, 8'h80, 8'h24, 8'h02, 8'h32,
			8'h02, 8'h24, 8'h02, 8'hFF, 8'hC8, 8'h84, 8'h02, 8'hFF, 8'h81, 8'h14, 8'h02, 8'h02, 8'h14, 8'h1A, 8'h14, 8'h02,
			8'h02, 8'h88, 8'h10, 8'h10, 8'h10, 8'h10, 8'h14, 8'h10, 8'h85, 8'h3C, 8'h81, 8'h44, 8'h85, 8'h4A, 8'h81, 8'h44,
			8'h88, 8'h28, 8'h24, 8'h20, 8'h46, 8'h42, 8'h40, 8'hC6, 8'h81, 8'h3C, 8'h02, 8'h02, 8'h44, 8'h02, 8'h02, 8'h02,
			8'h4A, 8'h02, 8'h46, 8'h36, 8'h36, 8'h38, 8'h38, 8'h02, 8'h3A, 8'h02, 8'h80, 8'h3C, 8'h3C, 8'h81, 8'h02, 8'h24,
			8'h02, 8'h02, 8'h2C, 8'h24, 8'h88, 8'h24, 8'h1E, 8'h46, 8'h36, 8'h38, 8'h3A, 8'hFF, 8'hC4, 8'h84, 8'h02, 8'hFF,
			8'hD8, 8'h81, 8'h06, 8'hFF, 8'hC6, 8'h88, 8'h06, 8'hFF, 8'hC7, 8'h81, 8'h06, 8'h06, 8'h80, 8'h06, 8'h06, 8'h81,
			8'h06, 8'h06, 8'h80, 8'h06, 8'h06, 8'h81, 8'h06, 8'h06, 8'hFF, 8'hC6, 8'h88, 8'h06, 8'hFF, 8'hE0, 8'h81, 8'h06,
			8'h06, 8'hFF, 8'h82, 8'h0F, 8'h81, 8'h06, 8'h06, 8'hEA, 8'h06, 8'h06, 8'h06, 8'h06, 8'hFF, 8'hC5, 8'h80, 8'h0E,
			8'h58, 8'hFF, 8'h00, 8'hC5, 8'h80, 8'h0E, 8'h58, 8'hFF, 8'h82, 8'h1C, 8'h1C, 8'hC3, 8'h82, 8'h1C, 8'h1C, 8'h81,
			8'h1C, 8'h1C, 8'h1C, 8'h02, 8'hFF, 8'hC7, 8'h88, 8'h1C, 8'hFF, 8'h00, 8'h83, 8'h02, 8'h80, 8'h0E, 8'h02, 8'h0E,
			8'h02, 8'h0C, 8'h02, 8'h0E, 8'h02, 8'h4E, 8'h02, 8'h02, 8'h02, 8'h0E, 8'h02, 8'h0C, 8'h02, 8'h02, 8'h02, 8'h0E,
			8'h02, 8'h0C, 8'h02, 8'h0E, 8'h02, 8'h4E, 8'h02, 8'h02, 8'h02, 8'h0E, 8'h02, 8'h0C, 8'h02, 8'h0E, 8'h02, 8'h0E,
			8'h02, 8'h0C, 8'h02, 8'h0E, 8'h02, 8'h4E, 8'h02, 8'h02, 8'h02, 8'h0E, 8'h02, 8'h0C, 8'h02, 8'h88, 8'h4E, 8'h18,
			8'h16, 8'h12, 8'h0E, 8'h0C, 8'h0E, 8'h83, 8'h02, 8'h81, 8'h3E, 8'h3E, 8'h82, 8'h46, 8'h1C, 8'h46, 8'h81, 8'h02,
			8'h38, 8'h3E, 8'h02, 8'h82, 8'h46, 8'h1C, 8'h82, 8'h48, 8'h48, 8'h81, 8'h3E, 8'h3E, 8'h82, 8'h38, 8'h88, 8'h24,
			8'h20, 8'h1C, 8'h48, 8'h46, 8'h42, 8'h3E, 8'h82, 8'h09, 8'h09, 8'hC6, 8'h82, 8'h03, 8'h0C, 8'hFF, 8'hC6, 8'h88,
			8'h06, 8'hFF, 8'hED, 8'h89, 8'h2A, 8'h02, 8'h04, 8'h0C, 8'h02, 8'h04, 8'h08, 8'h02, 8'h30, 8'h26, 8'h02, 8'h30,
			8'hFF, 8'h80, 8'h02, 8'hED, 8'h89, 8'h0C, 8'h02, 8'h12, 8'h4E, 8'h02, 8'h12, 8'h18, 8'h02, 8'h0E, 8'h08, 8'h02,
			8'h0E, 8'hFF, 8'h80, 8'h42, 8'h02, 8'h48, 8'h02, 8'h1E, 8'h02, 8'h24, 8'h02, 8'h02, 8'h02, 8'h2A, 8'h02, 8'hC6,
			8'h8C, 8'h30, 8'h2A, 8'hFF, 8'h00, 8'h80, 8'h24, 8'h02, 8'h2A, 8'h02, 8'h30, 8'h02, 8'h06, 8'h02, 8'h02, 8'h02,
			8'h0C, 8'h02, 8'hC6, 8'h8C, 8'h12, 8'h18, 8'hFF, 8'h80, 8'h56, 8'h54, 8'h52, 8'h50, 8'h81, 8'h02, 8'h80, 8'h5E,
			8'h5A, 8'h54, 8'h50, 8'h18, 8'h14, 8'h10, 8'h0A, 8'h06, 8'h30, 8'h2C, 8'h28, 8'h02, 8'h00, 8'h80, 8'h1A, 8'h18,
			8'h16, 8'h14, 8'h81, 8'h02, 8'h80, 8'h02, 8'h5E, 8'h5A, 8'h54, 8'h50, 8'h18, 8'h14, 8'h10, 8'h0A, 8'h06, 8'h30,
			8'h2C, 8'h28, 8'h82, 8'h1C, 8'h02, 8'h1C, 8'h02, 8'h02, 8'h1C, 8'h1C, 8'h00, 8'h81, 8'h10, 8'h0A, 8'h32, 8'h28,
			8'h80, 8'h32, 8'h02, 8'h32, 8'h02, 8'h82, 8'h32, 8'h81, 8'h06, 8'h02, 8'h06, 8'h02, 8'h82, 8'h32, 8'h81, 8'h54,
			8'h1A, 8'h10, 8'h0A, 8'h80, 8'h10, 8'h02, 8'h10, 8'h02, 8'h82, 8'h10, 8'h81, 8'h16, 8'h02, 8'h16, 8'h02, 8'h82,
			8'h0A, 8'h83, 8'h03, 8'h0C, 8'h82, 8'h03, 8'h0C, 8'h0C, 8'hC2, 8'h88, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C,
			8'h83, 8'h1C, 8'h80, 8'h04, 8'h04, 8'h2A, 8'h02, 8'h82, 8'h1C, 8'hFF, 8'h81, 8'h4C, 8'h02, 8'h4C, 8'h02, 8'h2A,
			8'h02, 8'h4C, 8'h1C, 8'h81, 8'h4C, 8'h02, 8'h4C, 8'h02, 8'h4C, 8'h00, 8'h88, 8'h2E, 8'h2E, 8'h2E, 8'h30, 8'h04,
			8'h30, 8'hC4, 8'h80, 8'h2E, 8'h04, 8'hFF, 8'h83, 8'h02, 8'h88, 8'h2E, 8'h2E, 8'h2E, 8'h30, 8'h04, 8'h30, 8'hC4,
			8'h80, 8'h2E, 8'h04, 8'hFF, 8'h83, 8'h02, 8'h84, 8'h02, 8'h02, 8'hC2, 8'h88, 8'h3E, 8'h3E, 8'h3E, 8'h42, 8'h46,
			8'h42, 8'h84, 8'h3E, 8'hFF, 8'h85, 8'h3E, 8'h81, 8'h3E, 8'h88, 8'h1C, 8'h46, 8'h1C, 8'h81, 8'h02, 8'h3E, 8'h3E,
			8'h3E, 8'h82, 8'h34, 8'h02, 8'hC2, 8'h88, 8'h06, 8'h06, 8'h06, 8'h06, 8'h06, 8'h06, 8'h82, 8'h06, 8'h06, 8'h06,
			8'h06, 8'hFF, 8'hC2, 8'h81, 8'h06, 8'h06, 8'h80, 8'h06, 8'h06, 8'h81, 8'h06, 8'h06, 8'h06, 8'h06, 8'h80, 8'h06,
			8'h06, 8'hFF, 8'h09, 8'h80, 8'h10, 8'h02, 8'h10, 8'h02, 8'h10, 8'h02, 8'h0C, 8'h0C, 8'h0C, 8'h02, 8'h0C, 8'h02,
			8'h14, 8'h14, 8'h14, 8'h02, 8'h14, 8'h02, 8'h85, 8'h10, 8'h00, 8'h80, 8'h32, 8'h02, 8'h32, 8'h02, 8'h32, 8'h02,
			8'hC2, 8'h32, 8'h32, 8'h32, 8'h02, 8'h32, 8'h02, 8'hFF, 8'h85, 8'h32, 8'h80, 8'h54, 8'h02, 8'h54, 8'h02, 8'h54,
			8'h02, 8'h50, 8'h50, 8'h50, 8'h02, 8'h50, 8'h02, 8'h56, 8'h56, 8'h56, 8'h02, 8'h56, 8'h02, 8'h85, 8'h54, 8'hC4,
			8'h85, 8'h0C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4C, 8'h58, 8'hF7, 8'h94, 8'hC0, 8'h00, 8'hC0, 8'hF7, 8'hC0
		};
		chr_bits = '{
			8'h1E, 8'h3F, 8'h7F, 8'h7F, 8'hFF, 8'hFF, 8'h7F, 8'h7F, 8'h00, 8'h00, 8'h02, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00,
			8'h3F, 8'h1E, 8'h04, 8'h02, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h00, 8'h00, 8'h04, 8'h02, 8'h07, 8'h0F, 8'h0F, 8'h0B,
			8'h1F, 8'h1F, 8'h07, 8'h03, 8'h01, 8'h01, 8'h00, 8'h00, 8'h1A, 8'h1E, 8'h07, 8'h00, 8'h00, 8'h04, 8'h07, 8'h03,
			8'h78, 8'h7C, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'h00, 8'h80, 8'h48, 8'h44, 8'h24, 8'h20, 8'h40, 8'h40,
			8'h7C, 8'h78, 8'h20, 8'h40, 8'h00, 8'h84, 8'h0C, 8'h0C, 8'h80, 8'h00, 8'h20, 8'h40, 8'hC0, 8'hE4, 8'hEC, 8'hEC,
			8'h06, 8'h20, 8'hC0, 8'h90, 8'hF0, 8'hF0, 8'hE0, 8'h00, 8'hFE, 8'hD8, 8'hB0, 8'h60, 8'h80, 8'h00, 8'h00, 8'h80,
			8'h7C, 8'h78, 8'h20, 8'h40, 8'h00, 8'h80, 8'h00, 8'h00, 8'h80, 8'h00, 8'h20, 8'h40, 8'hC0, 8'hE0, 8'hE0, 8'hE0,
			8'h00, 8'h26, 8'hC7, 8'h94, 8'hF0, 8'hF0, 8'hE0, 8'h00, 8'hE0, 8'hDE, 8'hBF, 8'h64, 8'h80, 8'h00, 8'h00, 8'h80,
			8'h00, 8'h00, 8'hE0, 8'h80, 8'hC0, 8'hE0, 8'hFC, 8'h0E, 8'hE0, 8'hC0, 8'h80, 8'h70, 8'hB8, 8'h18, 8'h1C, 8'h8E,
			8'h00, 8'h1E, 8'h3F, 8'h7F, 8'h7F, 8'hFF, 8'hFF, 8'h7F, 8'h00, 8'h00, 8'h00, 8'h02, 8'h01, 8'h01, 8'h00, 8'h00,
			8'h7F, 8'h3F, 8'h1E, 8'h04, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h04, 8'h07, 8'h0F, 8'h0F, 8'h0B,
			8'h78, 8'hFC, 8'h7E, 8'hBE, 8'hBF, 8'hDF, 8'hDE, 8'hBE, 8'h00, 8'h00, 8'h88, 8'h44, 8'h44, 8'h20, 8'h20, 8'h40,
			8'hBC, 8'h78, 8'h20, 8'h40, 8'h00, 8'h84, 8'h0C, 8'h0C, 8'h40, 8'h00, 8'h20, 8'h40, 8'hC0, 8'hE4, 8'hEC, 8'hEC,
			8'h00, 8'h78, 8'hBC, 8'hBE, 8'hDE, 8'hDF, 8'hBF, 8'hBE, 8'h00, 8'h00, 8'h40, 8'h48, 8'h24, 8'h24, 8'h40, 8'h40,
			8'h7E, 8'hFC, 8'h78, 8'h20, 8'h00, 8'h84, 8'h0C, 8'h0C, 8'h80, 8'h00, 8'h00, 8'h20, 8'hC0, 8'hE4, 8'hEC, 8'hEC,
			8'h03, 8'h07, 8'h0F, 8'h0F, 8'h1F, 8'h1F, 8'h0F, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h07, 8'h03, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h00, 8'h00, 8'h01, 8'h01, 8'h07, 8'h0F, 8'h0F, 8'h0B,
			8'hC0, 8'hE0, 8'hF0, 8'hF0, 8'hF8, 8'hF8, 8'hF0, 8'hF0, 8'h00, 8'h00, 8'h40, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00,
			8'hE0, 8'hC0, 8'h00, 8'h00, 8'h00, 8'h84, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE4, 8'hEC, 8'hEC,
			8'h00, 8'h01, 8'h03, 8'h07, 8'h07, 8'h0F, 8'h0F, 8'h07, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h07, 8'h03, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h01, 8'h07, 8'h0F, 8'h0F, 8'h0B,
			8'h00, 8'hE0, 8'hF0, 8'hF8, 8'hF8, 8'hFC, 8'hFC, 8'hF8, 8'h00, 8'h00, 8'h00, 8'h20, 8'h10, 8'h10, 8'h00, 8'h00,
			8'hF8, 8'hF0, 8'hE0, 8'h00, 8'h00, 8'h84, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE4, 8'hEC, 8'hEC,
			8'h1F, 8'h0F, 8'h07, 8'h01, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h01, 8'h07, 8'h0F, 8'h0F, 8'h0B,
			8'hE0, 8'hC0, 8'h80, 8'h00, 8'h00, 8'h84, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE4, 8'hEC, 8'hEC,
			8'hE0, 8'hC0, 8'h00, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE0, 8'hE0, 8'hE0,
			8'h07, 8'h0F, 8'h1F, 8'h1F, 8'h3F, 8'h3F, 8'h1F, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h0F, 8'h05, 8'h00, 8'h02, 8'h00, 8'h3C, 8'h7C, 8'h7C, 8'h00, 8'h00, 8'h1F, 8'h3F, 8'h3F, 8'h2B, 8'h6B, 8'h7B,
			8'h1E, 8'h6E, 8'h5C, 8'h1F, 8'h3F, 8'h1F, 8'h03, 8'h00, 8'h1E, 8'h61, 8'h63, 8'h84, 8'hC0, 8'h60, 8'h20, 8'h01,
			8'h80, 8'hD8, 8'hEC, 8'hEE, 8'hF6, 8'hF7, 8'hEF, 8'hEE, 8'h00, 8'h20, 8'h90, 8'h58, 8'h4C, 8'h0C, 8'h10, 8'h10,
			8'hDE, 8'hBC, 8'h78, 8'h10, 8'h20, 8'h40, 8'h00, 8'h00, 8'h20, 8'h40, 8'h00, 8'h90, 8'hA0, 8'hC0, 8'h80, 8'h00,
			8'h60, 8'h60, 8'h40, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'hE0, 8'hE0, 8'h40, 8'h00, 8'h00, 8'h40, 8'hC0, 8'h80,
			8'h3C, 8'h18, 8'h1C, 8'h7C, 8'h7D, 8'h3F, 8'h06, 8'h00, 8'h3C, 8'h06, 8'h23, 8'h47, 8'h4E, 8'h00, 8'h70, 8'h0E,
			8'h0F, 8'h07, 8'h02, 8'h00, 8'h02, 8'h00, 8'h3C, 8'h7C, 8'h00, 8'h00, 8'h02, 8'h1F, 8'h3F, 8'h3F, 8'h2B, 8'h6B,
			8'h7C, 8'h1E, 8'h6D, 8'h61, 8'h03, 8'h1F, 8'h0D, 8'h00, 8'h7B, 8'h1E, 8'h62, 8'h7E, 8'h3C, 8'h00, 8'h00, 8'h1C,
			8'hDE, 8'hBC, 8'h78, 8'h10, 8'h20, 8'h40, 8'h00, 8'h00, 8'h20, 8'h40, 8'h00, 8'h10, 8'hA0, 8'hC0, 8'h80, 8'h80,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'h80, 8'h80, 8'h00, 8'h00, 8'h00, 8'h80, 8'h80, 8'h40, 8'h60, 8'h20, 8'h00,
			8'h1E, 8'h3F, 8'h7F, 8'h7F, 8'hFF, 8'hFF, 8'h7F, 8'h7F, 8'h00, 8'h00, 8'h02, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00,
			8'h3F, 8'h1E, 8'h01, 8'h00, 8'h01, 8'h00, 8'h1E, 8'h3E, 8'h00, 8'h01, 8'h01, 8'h0F, 8'h1F, 8'h1F, 8'h15, 8'h35,
			8'h3E, 8'h0F, 8'h36, 8'h2F, 8'h1F, 8'h1F, 8'h0F, 8'h08, 8'h3D, 8'h0F, 8'h31, 8'h30, 8'h44, 8'h60, 8'h70, 8'h30,
			8'h00, 8'h60, 8'hB0, 8'hB8, 8'hD8, 8'hDC, 8'hBC, 8'hB8, 8'h00, 8'h80, 8'h40, 8'h60, 8'h30, 8'h30, 8'h40, 8'h40,
			8'h78, 8'hF0, 8'hE0, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'hA0, 8'hC0, 8'hC0, 8'hC0, 8'hC0,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'hE0, 8'h40, 8'h00, 8'h80, 8'h00, 8'hC0, 8'hE0, 8'h60, 8'hE0, 8'h40, 8'h00,
			8'h1F, 8'h07, 8'h0E, 8'h1C, 8'h18, 8'h1C, 8'h08, 8'h00, 8'h1E, 8'h07, 8'h01, 8'h03, 8'h07, 8'h1F, 8'h0B, 8'h00,
			8'hC0, 8'h80, 8'h30, 8'h10, 8'h88, 8'h18, 8'h38, 8'h30, 8'h00, 8'h80, 8'hB0, 8'hF0, 8'hE0, 8'hE0, 8'hC0, 8'h40,
			8'h01, 8'h00, 8'h00, 8'h02, 8'h00, 8'h3C, 8'h7C, 8'h7C, 8'h00, 8'h00, 8'h1F, 8'h3F, 8'h3F, 8'h2B, 8'h6B, 8'h7B,
			8'hFE, 8'hFC, 8'h78, 8'h10, 8'h20, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h90, 8'hA0, 8'hC0, 8'h80, 8'h00,
			8'h01, 8'h00, 8'h00, 8'h00, 8'h02, 8'h00, 8'h3C, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h1F, 8'h3F, 8'h3F, 8'h2B, 8'h6B,
			8'hFE, 8'hFC, 8'h78, 8'h10, 8'h20, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'hA0, 8'hC0, 8'h80, 8'h80,
			8'h3F, 8'h1E, 8'h01, 8'h00, 8'h01, 8'h00, 8'h1E, 8'h3E, 8'h00, 8'h00, 8'h01, 8'h0F, 8'h1F, 8'h1F, 8'h15, 8'h35,
			8'h00, 8'h00, 8'h80, 8'h80, 8'hC0, 8'hC0, 8'h80, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'hC0, 8'hC0, 8'hC0, 8'hC0,
			8'h3F, 8'h1E, 8'h04, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h1F, 8'h00, 8'h00, 8'h04, 8'h07, 8'h0F, 8'h0F, 8'h0A, 8'h1A,
			8'h1F, 8'h07, 8'h03, 8'h07, 8'h1F, 8'h1F, 8'h0E, 8'h00, 8'h1E, 8'h07, 8'h0C, 8'h18, 8'h1A, 8'h10, 8'h00, 8'h1C,
			8'h7C, 8'h78, 8'h40, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h80, 8'h00, 8'h40, 8'hC0, 8'hE0, 8'hE0, 8'hE0, 8'hE0,
			8'h00, 8'h80, 8'h00, 8'h80, 8'h80, 8'hE0, 8'hE0, 8'h00, 8'hC0, 8'h80, 8'hC0, 8'h60, 8'hE0, 8'hC0, 8'h00, 8'h70,
			8'h3F, 8'h1E, 8'h04, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h1F, 8'h00, 8'h00, 8'h04, 8'h07, 8'h0F, 8'h0F, 8'h0A, 8'h1A,
			8'h7E, 8'hFC, 8'h78, 8'h20, 8'h80, 8'h00, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'hE0,
			8'h7F, 8'h3F, 8'h1E, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h0A, 8'h1A,
			8'hBC, 8'h78, 8'h40, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h40, 8'h00, 8'h40, 8'hC0, 8'hE0, 8'hE0, 8'hE0, 8'hE0,
			8'h07, 8'h03, 8'h01, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h0A, 8'h1A,
			8'hF8, 8'hF0, 8'hE0, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE0, 8'hE0, 8'hE0, 8'hE0,
			8'h1F, 8'h0F, 8'h07, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h0A, 8'h1A,
			8'hE0, 8'hC0, 8'h80, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE0, 8'hE0, 8'hE0, 8'hE0,
			8'h07, 8'h03, 8'h01, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h1F, 8'h00, 8'h00, 8'h01, 8'h07, 8'h0F, 8'h0F, 8'h0A, 8'h1A,
			8'hE0, 8'hC0, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE0, 8'hE0, 8'hE0, 8'hE0,
			8'hCF, 8'h4F, 8'h07, 8'h0F, 8'h07, 8'h07, 8'h03, 8'h00, 8'hF5, 8'h77, 8'h1F, 8'h03, 8'h1C, 8'h18, 8'h0C, 8'h04,
			8'hE6, 8'hE4, 8'hC0, 8'hE0, 8'hC0, 8'hC0, 8'h80, 8'h00, 8'h5E, 8'hDC, 8'hF0, 8'h80, 8'h70, 8'h30, 8'h60, 8'h40,
			8'h0F, 8'h0F, 8'h07, 8'hEF, 8'h27, 8'h07, 8'h03, 8'h00, 8'h05, 8'h37, 8'h7F, 8'hE3, 8'h3C, 8'h18, 8'h0C, 8'h04,
			8'hE0, 8'hE0, 8'hC0, 8'hEE, 8'hC8, 8'hC0, 8'h80, 8'h00, 8'h40, 8'hD8, 8'hFC, 8'h8E, 8'h78, 8'h30, 8'h60, 8'h40,
			8'h0F, 8'h07, 8'h03, 8'h07, 8'h1F, 8'h37, 8'h03, 8'h00, 8'h07, 8'h0F, 8'h1F, 8'h1C, 8'h18, 8'h38, 8'h0C, 8'h04,
			8'hE0, 8'hC0, 8'h80, 8'hC0, 8'hF0, 8'hD8, 8'h80, 8'h00, 8'hC0, 8'hE0, 8'hF0, 8'h70, 8'h30, 8'h38, 8'h60, 8'h40,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h05,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h40, 8'h00, 8'hE0, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE0, 8'hE0, 8'h40,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h05, 8'h07,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h40, 8'h00, 8'hE0, 8'hE0, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hA0, 8'hE0, 8'h40, 8'hC0,
			8'h0B, 8'hDA, 8'hE0, 8'h6D, 8'h29, 8'h03, 8'h5B, 8'hC5, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h78, 8'hFC, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h08, 8'h04, 8'h04, 8'h00, 8'h00,
			8'h03, 8'h07, 8'h0F, 8'h0F, 8'h1F, 8'h1F, 8'h0F, 8'h0F, 8'h03, 8'h07, 8'h0F, 8'h0F, 8'h1F, 8'h1F, 8'h0F, 8'h0F,
			8'h07, 8'h03, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h37, 8'h07, 8'h03, 8'h01, 8'h01, 8'h00, 8'h00, 8'h0E, 8'h0C,
			8'hFF, 8'h1F, 8'h07, 8'h00, 8'h00, 8'h04, 8'h07, 8'h03, 8'h01, 8'h1F, 8'h07, 8'h03, 8'h01, 8'h01, 8'h00, 8'h00,
			8'hC0, 8'hE0, 8'hB0, 8'hD0, 8'hD8, 8'hF8, 8'hF0, 8'hF0, 8'hC0, 8'hE0, 8'hF0, 8'hF0, 8'hF8, 8'hF8, 8'hF0, 8'hF0,
			8'hE0, 8'hC0, 8'h00, 8'h00, 8'h80, 8'h84, 8'h2C, 8'hEC, 8'hE0, 8'hC0, 8'h00, 8'h20, 8'h20, 8'h60, 8'hC0, 8'h00,
			8'hDE, 8'hD8, 8'hB0, 8'h60, 8'h00, 8'h00, 8'h00, 8'h80, 8'hD8, 8'hF8, 8'hF0, 8'hF0, 8'hF0, 8'hF0, 8'hE0, 8'h00,
			8'h01, 8'h03, 8'h07, 8'h07, 8'h0F, 8'h0F, 8'h07, 8'h07, 8'h01, 8'h03, 8'h07, 8'h07, 8'h0F, 8'h0F, 8'h07, 8'h07,
			8'h03, 8'h01, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h37, 8'h03, 8'h01, 8'h00, 8'h01, 8'h00, 8'h00, 8'h0E, 8'h0C,
			8'hE0, 8'hF0, 8'hD8, 8'hE8, 8'hEC, 8'hFC, 8'hF8, 8'hF8, 8'hE0, 8'hF0, 8'hF8, 8'hF8, 8'hFC, 8'hFC, 8'hF8, 8'hF8,
			8'hF0, 8'hE0, 8'h00, 8'h00, 8'h80, 8'h84, 8'h2C, 8'hEC, 8'hF0, 8'hE0, 8'h80, 8'h20, 8'h20, 8'h60, 8'hC0, 8'h00,
			8'hC0, 8'hDE, 8'hBF, 8'h64, 8'h00, 8'h00, 8'h00, 8'h80, 8'hC0, 8'hF8, 8'hF8, 8'hF0, 8'hF0, 8'hF0, 8'hE0, 8'h00,
			8'h00, 8'h07, 8'h0F, 8'h1F, 8'h1F, 8'h3F, 8'h3F, 8'h1F, 8'h00, 8'h07, 8'h0F, 8'h1F, 8'h1F, 8'h3F, 8'h3F, 8'h1F,
			8'h1F, 8'h0F, 8'h07, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h37, 8'h1F, 8'h0F, 8'h07, 8'h01, 8'h00, 8'h00, 8'h0E, 8'h0C,
			8'h00, 8'h80, 8'hC0, 8'h60, 8'hA0, 8'hB0, 8'hF0, 8'hE0, 8'h00, 8'h80, 8'hC0, 8'hE0, 8'hE0, 8'hF0, 8'hF0, 8'hE0,
			8'hE0, 8'hC0, 8'h80, 8'h00, 8'h80, 8'h84, 8'h2C, 8'hEC, 8'hE0, 8'hC0, 8'h80, 8'h20, 8'h20, 8'h60, 8'hC0, 8'h00,
			8'hC0, 8'hC0, 8'h80, 8'h60, 8'h32, 8'h1E, 8'h1C, 8'h88, 8'hC0, 8'hC0, 8'hE0, 8'hF0, 8'hF8, 8'hF8, 8'hF0, 8'h00,
			8'hE0, 8'hC0, 8'h00, 8'h00, 8'h80, 8'h80, 8'h20, 8'hE0, 8'hE0, 8'hC0, 8'h00, 8'h20, 8'h20, 8'h60, 8'hC0, 8'h00,
			8'h02, 8'h0E, 8'h0B, 8'h00, 8'h01, 8'h07, 8'h0F, 8'h0F, 8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h0E,
			8'h3B, 8'h7F, 8'h5F, 8'h46, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h01, 8'h1F, 8'h07, 8'h01, 8'h00, 8'h00, 8'h00,
			8'hC0, 8'hA0, 8'h40, 8'h80, 8'h00, 8'h80, 8'h80, 8'h20, 8'h00, 8'h40, 8'h80, 8'h80, 8'h00, 8'h20, 8'h60, 8'hD8,
			8'h60, 8'h80, 8'h60, 8'hE0, 8'hD8, 8'hDC, 8'hCC, 8'h60, 8'h9C, 8'hFE, 8'hFE, 8'hFE, 8'hE6, 8'hE0, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h28, 8'h54, 8'hD4, 8'hBA, 8'hBB, 8'h7D, 8'h00, 8'h00, 8'h10, 8'h28, 8'h28, 8'h44, 8'h44, 8'h02,
			8'h01, 8'h00, 8'h00, 8'h01, 8'h01, 8'h07, 8'h0F, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h00, 8'h00, 8'h0E,
			8'h50, 8'hB0, 8'h80, 8'h00, 8'h00, 8'h80, 8'h80, 8'h20, 8'hA0, 8'h80, 8'h80, 8'h00, 8'h00, 8'h20, 8'h60, 8'hD8,
			8'h06, 8'h1D, 8'h3B, 8'h7B, 8'h77, 8'hF7, 8'hF7, 8'hE3, 8'h01, 8'h02, 8'h04, 8'h04, 8'h08, 8'h08, 8'h00, 8'h00,
			8'h81, 8'h41, 8'h21, 8'h11, 8'h09, 8'h07, 8'h0F, 8'h0F, 8'h00, 8'h41, 8'h21, 8'h11, 8'h09, 8'h00, 8'h00, 8'h0E,
			8'hC0, 8'h70, 8'hB8, 8'hBC, 8'hDC, 8'hDE, 8'hDE, 8'h8E, 8'h00, 8'h80, 8'h40, 8'h40, 8'h20, 8'h20, 8'h00, 8'h00,
			8'h02, 8'h04, 8'h08, 8'h10, 8'h00, 8'h80, 8'h80, 8'h20, 8'h00, 8'h04, 8'h08, 8'h10, 8'h20, 8'h20, 8'h60, 8'hD8,
			8'h0C, 8'h06, 8'h43, 8'h63, 8'h67, 8'hE7, 8'hF7, 8'hE3, 8'h02, 8'h81, 8'h20, 8'h10, 8'h10, 8'h18, 8'h00, 8'h00,
			8'h18, 8'h30, 8'h31, 8'h73, 8'h76, 8'hE6, 8'hFF, 8'h8F, 8'h00, 8'h04, 8'h82, 8'h84, 8'h88, 8'h18, 8'h00, 8'h00,
			8'h10, 8'h18, 8'h0F, 8'h07, 8'h33, 8'h23, 8'h63, 8'h61, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h02, 8'h1B, 8'h19,
			8'h41, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h1F, 8'h1F, 8'h0F, 8'h0F, 8'h07, 8'h00, 8'h00,
			8'h00, 8'hE0, 8'hF0, 8'h78, 8'hF8, 8'hE0, 8'hF0, 8'hF8, 8'h00, 8'h00, 8'hC0, 8'hC0, 8'hC2, 8'h1A, 8'hCE, 8'hE0,
			8'hE0, 8'h00, 8'h60, 8'hF0, 8'h38, 8'h38, 8'h10, 8'h00, 8'hE0, 8'hC0, 8'hE0, 8'hF0, 8'hB0, 8'h00, 8'h00, 8'h00,
			8'hE4, 8'h0C, 8'h3E, 8'hF8, 8'h60, 8'h00, 8'h00, 8'h00, 8'hE0, 8'hC0, 8'hF8, 8'hF8, 8'hE0, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h0F, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01,
			8'h00, 8'h00, 8'h78, 8'hF8, 8'hF2, 8'h76, 8'hFC, 8'hFC, 8'h00, 8'h02, 8'h02, 8'h06, 8'hEC, 8'hC8, 8'h1C, 8'hFC,
			8'h60, 8'h18, 8'h38, 8'h30, 8'h70, 8'hE0, 8'hC6, 8'h1C, 8'h7E, 8'h3E, 8'h3F, 8'h3F, 8'h7F, 8'h1F, 8'hC8, 8'hE0,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h0F, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h00,
			8'h00, 8'h78, 8'hF8, 8'hF2, 8'h76, 8'hFC, 8'hF0, 8'h6C, 8'h02, 8'h02, 8'h06, 8'hEC, 8'hC8, 8'h1C, 8'hFE, 8'h7E,
			8'hFC, 8'hD8, 8'h40, 8'h40, 8'h40, 8'hC2, 8'hC6, 8'h0C, 8'h1F, 8'h7F, 8'h3F, 8'h3F, 8'h1F, 8'hCC, 8'hC0, 8'hE0,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h1E, 8'h1E, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h1E, 8'h1E, 8'h0D,
			8'h00, 8'h00, 8'h1C, 8'h3A, 8'h3A, 8'h3E, 8'h3E, 8'h1C, 8'h00, 8'h00, 8'h1C, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h1D,
			8'h3C, 8'h76, 8'h7A, 8'hFB, 8'hFF, 8'h7E, 8'h7E, 8'h3C, 8'h3C, 8'h7E, 8'h7E, 8'hFF, 8'hFF, 8'h7E, 8'h7E, 8'h3D,
			8'h00, 8'h00, 8'h08, 8'h38, 8'h50, 8'h72, 8'hE3, 8'hE7, 8'h00, 8'h00, 8'h06, 8'h06, 8'h2E, 8'h0C, 8'h1C, 8'h18,
			8'h0B, 8'h1E, 8'h3F, 8'h7F, 8'h7E, 8'hFC, 8'hFC, 8'hFD, 8'h0C, 8'h0D, 8'h00, 8'h00, 8'h01, 8'h03, 8'h2B, 8'h13,
			8'h80, 8'hC0, 8'h80, 8'h10, 8'h20, 8'h40, 8'h80, 8'h00, 8'h00, 8'h30, 8'h70, 8'hF0, 8'hF8, 8'hF8, 8'hF0, 8'hE0,
			8'h00, 8'h0F, 8'h3D, 8'h3F, 8'h76, 8'h76, 8'hFC, 8'hFC, 8'h00, 8'h00, 8'h02, 8'h00, 8'h39, 8'h39, 8'h3B, 8'h03,
			8'hFC, 8'hFC, 8'hFC, 8'hFE, 8'hFF, 8'h7F, 8'h7F, 8'h3F, 8'h03, 8'h03, 8'h03, 8'h09, 8'h08, 8'h04, 8'h04, 8'h08,
			8'h00, 8'h90, 8'h00, 8'h20, 8'h00, 8'h40, 8'h00, 8'h84, 8'h60, 8'h70, 8'hE0, 8'hE0, 8'hC0, 8'hC0, 8'h80, 8'h84,
			8'h10, 8'h40, 8'h00, 8'h18, 8'hFC, 8'hAC, 8'hAC, 8'hAC, 8'h1E, 8'h7E, 8'hFC, 8'hE0, 8'h00, 8'h50, 8'h50, 8'h50,
			8'h00, 8'h07, 8'h1D, 8'h3E, 8'h6E, 8'h7E, 8'hFE, 8'hFC, 8'h00, 8'h00, 8'h02, 8'h31, 8'h79, 8'h79, 8'h79, 8'h33,
			8'hFC, 8'hF8, 8'hF8, 8'hF0, 8'hF8, 8'hFC, 8'hFF, 8'h7F, 8'h03, 8'h07, 8'h06, 8'h0E, 8'h17, 8'h13, 8'h20, 8'h00,
			8'h79, 8'h71, 8'h21, 8'h13, 8'h73, 8'h07, 8'h07, 8'h01, 8'h06, 8'h0E, 8'h1E, 8'hFC, 8'hFC, 8'hF8, 8'h78, 8'h70,
			8'h00, 8'h20, 8'h00, 8'h20, 8'h00, 8'h40, 8'h00, 8'h40, 8'hC0, 8'hE0, 8'hC0, 8'hE0, 8'hC0, 8'hC0, 8'h80, 8'hC0,
			8'h00, 8'h00, 8'h02, 8'hA8, 8'h00, 8'h00, 8'hF8, 8'hFC, 8'h00, 8'h00, 8'h02, 8'hAF, 8'hFF, 8'hFE, 8'h00, 8'h00,
			8'hFC, 8'hF6, 8'hD6, 8'hDB, 8'hEB, 8'hEB, 8'hEB, 8'hEA, 8'h00, 8'h08, 8'h28, 8'h24, 8'h14, 8'h14, 8'h14, 8'h14,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h0F, 8'h1F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h3F, 8'h7F, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'h01, 8'h01, 8'h01, 8'h00, 8'h02, 8'h04, 8'h05, 8'h09,
			8'h00, 8'h00, 8'h00, 8'h00, 8'hE0, 8'hF0, 8'hF8, 8'hFC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0,
			8'hFC, 8'hBE, 8'hBA, 8'hFE, 8'h80, 8'h00, 8'h00, 8'h55, 8'hE0, 8'hE0, 8'hE4, 8'hC0, 8'h7E, 8'hFF, 8'hFF, 8'hD5,
			8'h00, 8'h20, 8'h20, 8'h10, 8'h10, 8'h1F, 8'h1F, 8'h0F, 8'h78, 8'h7C, 8'hFC, 8'hFC, 8'h78, 8'h60, 8'h20, 8'h00,
			8'h0F, 8'h07, 8'h07, 8'h07, 8'h0C, 8'h0C, 8'h0C, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h03, 8'h03, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hF0, 8'hF8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60,
			8'hFC, 8'hFC, 8'hFE, 8'hFE, 8'h7F, 8'hBF, 8'h3F, 8'h3F, 8'h10, 8'h10, 8'h08, 8'h08, 8'h80, 8'hC0, 8'hC0, 8'hC0,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h10, 8'h10, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hFE, 8'hFE, 8'h7C, 8'h38,
			8'h10, 8'h38, 8'h38, 8'h78, 8'h7C, 8'h7C, 8'h7E, 8'h7F, 8'h00, 8'h00, 8'h00, 8'h10, 8'h10, 8'h08, 8'h00, 8'h00,
			8'h03, 8'h07, 8'h06, 8'h04, 8'h0C, 8'h08, 8'h00, 8'h00, 8'h03, 8'h07, 8'h06, 8'h04, 8'h0C, 8'h08, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h07, 8'h06, 8'h04, 8'h0C, 8'h08, 8'h00, 8'h00,
			8'h03, 8'h07, 8'h06, 8'h0E, 8'h0C, 8'h1C, 8'h18, 8'h38, 8'h03, 8'h07, 8'h06, 8'h0E, 8'h0C, 8'h1C, 8'h18, 8'h38,
			8'h3C, 8'h0E, 8'h03, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h0E, 8'h03, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h07, 8'h06, 8'h0E, 8'h0C, 8'h1C, 8'h18, 8'h38,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h0E, 8'h03, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h03, 8'h07, 8'h06, 8'h0E, 8'h0C, 8'h1C, 8'h18, 8'h38, 8'h03, 8'h07, 8'h06, 8'h0E, 8'h0C, 8'h1C, 8'h18, 8'h38,
			8'h3C, 8'h0F, 8'h03, 8'h06, 8'h06, 8'h0C, 8'h0C, 8'h18, 8'h3C, 8'h0F, 8'h03, 8'h06, 8'h06, 8'h0C, 8'h0C, 8'h18,
			8'h18, 8'h30, 8'h30, 8'h20, 8'h60, 8'h40, 8'hC0, 8'h80, 8'h18, 8'h30, 8'h30, 8'h20, 8'h60, 8'h40, 8'hC0, 8'h80,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h07, 8'h06, 8'h0E, 8'h0C, 8'h1C, 8'h18, 8'h38,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h0F, 8'h03, 8'h06, 8'h06, 8'h0C, 8'h0C, 8'h18,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h30, 8'h30, 8'h20, 8'h60, 8'h40, 8'hC0, 8'h80,
			8'h00, 8'h00, 8'h10, 8'h1C, 8'h38, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h3C, 8'h18, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h18, 8'h3E, 8'h7C, 8'h18, 8'h08, 8'h00,
			8'h52, 8'h11, 8'h98, 8'h3F, 8'hFC, 8'h19, 8'h88, 8'h4A, 8'h52, 8'h19, 8'hBC, 8'h7F, 8'hFE, 8'h3D, 8'h98, 8'h4A,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h42, 8'h2C, 8'h38, 8'h1C, 8'h34, 8'h42, 8'h00,
			8'h81, 8'h66, 8'h7E, 8'h3C, 8'h3C, 8'h7E, 8'h66, 8'h81, 8'h81, 8'h66, 8'h7E, 8'h3C, 8'h3C, 8'h7E, 8'h66, 8'h81,
			8'h00, 8'h00, 8'h00, 8'h0F, 8'hCF, 8'h4F, 8'h07, 8'h0F, 8'h07, 8'h0F, 8'h0F, 8'h05, 8'hF5, 8'h77, 8'h1F, 8'h03,
			8'h00, 8'h40, 8'h00, 8'hE0, 8'hE6, 8'hE4, 8'hC0, 8'hE0, 8'hC0, 8'hE0, 8'hE0, 8'h40, 8'h5E, 8'hDC, 8'hF0, 8'h80,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0D, 8'h0D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F,
			8'h16, 8'h33, 8'h12, 8'h09, 8'h06, 8'h01, 8'h0B, 8'h04, 8'h17, 8'h33, 8'h12, 8'h09, 8'h06, 8'h01, 8'h0B, 8'h04,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'h60, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hE0, 8'hE0,
			8'hD0, 8'h98, 8'h90, 8'h20, 8'hC0, 8'h00, 8'hA0, 8'h40, 8'hD0, 8'h98, 8'h90, 8'h20, 8'hC0, 8'h00, 8'hA0, 8'h40,
			8'h03, 8'h07, 8'h0F, 8'h0F, 8'h1F, 8'h1F, 8'h1F, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC0, 8'hE0, 8'hB0, 8'h90, 8'hD8, 8'hD8, 8'hF8, 8'hF8, 8'h00, 8'h00, 8'h40, 8'h60, 8'h20, 8'h20, 8'h00, 8'h00,
			8'hFF, 8'hFF, 8'h7E, 8'h3C, 8'h10, 8'h08, 8'h04, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h08, 8'h04, 8'h04,
			8'hFF, 8'hFF, 8'h7E, 8'h3C, 8'h10, 8'h10, 8'h08, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h10, 8'h08, 8'h08,
			8'h04, 8'h06, 8'h32, 8'h3A, 8'h18, 8'h02, 8'h63, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h18, 8'h11, 8'h04, 8'h4C, 8'h1C, 8'h18, 8'h0A, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h04, 8'h66, 8'h4A, 8'h18, 8'h10, 8'h48, 8'h40, 8'h00, 8'h04, 8'h6E, 8'h7E, 8'h3C, 8'h3C, 8'h7C, 8'h6E, 8'hEF,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h66, 8'hC8, 8'h92, 8'h84, 8'h00, 8'h00, 8'h00, 8'h00, 8'h66, 8'hEE, 8'hFF, 8'hFF,
			8'h10, 8'h10, 8'h08, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7E, 8'h7C, 8'h3C, 8'h3C, 8'h2C, 8'h2C, 8'h2C, 8'h2C,
			8'h00, 8'h03, 8'h07, 8'h04, 8'h00, 8'h02, 8'h00, 8'h00, 8'h00, 8'h03, 8'h07, 8'h07, 8'h07, 8'h03, 8'h01, 8'h00,
			8'h0C, 8'h1A, 8'h90, 8'h90, 8'hA6, 8'h4D, 8'h48, 8'h45, 8'h0C, 8'h1E, 8'h9E, 8'h9C, 8'hBE, 8'hFF, 8'hFF, 8'hFF,
			8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hF8, 8'h70, 8'h70, 8'h30, 8'h20, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h3A, 8'h10,
			8'h00, 8'h00, 8'h40, 8'h80, 8'h80, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h78, 8'hF4, 8'hE0, 8'h60, 8'h00, 8'h00,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h0B,
			8'hFE, 8'hFC, 8'h78, 8'h20, 8'h00, 8'h84, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h20, 8'hC0, 8'hE4, 8'hEC, 8'hEC,
			8'h1E, 8'h3F, 8'h7F, 8'h7F, 8'hFF, 8'hFF, 8'h7F, 8'h7F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h3F, 8'h1E, 8'h04, 8'h07, 8'h0F, 8'h0F, 8'h0F, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h1F, 8'h07, 8'h0F, 8'h1F, 8'h1F, 8'h1F, 8'h0E, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h78, 8'hFC, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFC, 8'h78, 8'h40, 8'hC0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC0, 8'h80, 8'hC0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'h70, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h03, 8'h07, 8'h0F, 8'h0F, 8'h1F, 8'h1F, 8'h0F, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h07, 8'h03, 8'h01, 8'h07, 8'h0F, 8'h0F, 8'h0F, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC0, 8'hE0, 8'hF0, 8'hF0, 8'hF8, 8'hF8, 8'hF0, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hE0, 8'hC0, 8'h00, 8'hC0, 8'hE0, 8'hE0, 8'hE0, 8'hE0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h0C, 8'h10, 8'h21, 8'h20, 8'h40, 8'h40, 8'h48,
			8'h00, 8'h00, 8'h00, 8'hC0, 8'hE0, 8'h70, 8'h30, 8'h30, 8'hC0, 8'h30, 8'h08, 8'hC4, 8'h24, 8'h12, 8'h12, 8'h12,
			8'h10, 8'h10, 8'h08, 8'h08, 8'h06, 8'h01, 8'h00, 8'h00, 8'h48, 8'h48, 8'h44, 8'h26, 8'h21, 8'h10, 8'h0C, 8'h03,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'h02, 8'h02, 8'h02, 8'h04, 8'hC4, 8'h08, 8'h30, 8'hC0,
			8'h00, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h26, 8'h72, 8'h10, 8'h00, 8'hC0, 8'h60, 8'h00,
			8'h00, 8'hFF, 8'h8B, 8'hB9, 8'h88, 8'hBA, 8'h8B, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'hFC, 8'h4C, 8'h54, 8'h54, 8'h54, 8'h4C, 8'hFC, 8'hFE, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02,
			8'h00, 8'hFE, 8'h88, 8'hA4, 8'h84, 8'hA4, 8'h88, 8'hFE, 8'hFF, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01,
			8'h00, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h18, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08,
			8'h3F, 8'h60, 8'h40, 8'h40, 8'h40, 8'h60, 8'h3F, 8'h00, 8'h3F, 8'h7F, 8'h60, 8'h60, 8'h60, 8'h7F, 8'h3F, 8'h00,
			8'hFC, 8'h06, 8'h02, 8'h02, 8'h02, 8'h06, 8'hFC, 8'h00, 8'hFC, 8'hFE, 8'h06, 8'h06, 8'h06, 8'hFE, 8'hFC, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h02, 8'h05, 8'h01, 8'h02, 8'h01, 8'h01, 8'h05, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h07, 8'h04, 8'h04, 8'h06, 8'h01, 8'h01, 8'h05, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h07, 8'h05, 8'h01, 8'h01, 8'h02, 8'h02, 8'h02, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h12, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h17, 8'h34, 8'h14, 8'h16, 8'h11, 8'h11, 8'h15, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h22, 8'h55, 8'h55, 8'h15, 8'h25, 8'h45, 8'h45, 8'h72, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h72, 8'h45, 8'h45, 8'h65, 8'h15, 8'h15, 8'h55, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h22, 8'h55, 8'h55, 8'h55, 8'h55, 8'h55, 8'h55, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'h38, 8'h4C, 8'hC6, 8'hC6, 8'hC6, 8'h64, 8'h38, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h18, 8'h38, 8'h18, 8'h18, 8'h18, 8'h18, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h7C, 8'hC6, 8'h0E, 8'h3C, 8'h78, 8'hE0, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h7E, 8'h0C, 8'h18, 8'h3C, 8'h06, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h1C, 8'h3C, 8'h6C, 8'hCC, 8'hFE, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFC, 8'hC0, 8'hFC, 8'h06, 8'h06, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h3C, 8'h60, 8'hC0, 8'hFC, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFE, 8'hC6, 8'h0C, 8'h18, 8'h30, 8'h30, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h78, 8'hC4, 8'hE4, 8'h78, 8'h86, 8'h86, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h7C, 8'hC6, 8'hC6, 8'h7E, 8'h06, 8'h0C, 8'h78, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h38, 8'h6C, 8'hC6, 8'hC6, 8'hFE, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFC, 8'hC6, 8'hC6, 8'hFC, 8'hC6, 8'hC6, 8'hFC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h3C, 8'h66, 8'hC0, 8'hC0, 8'hC0, 8'h66, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hF8, 8'hCC, 8'hC6, 8'hC6, 8'hC6, 8'hCC, 8'hF8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFE, 8'hC0, 8'hC0, 8'hFC, 8'hC0, 8'hC0, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFE, 8'hC0, 8'hC0, 8'hFC, 8'hC0, 8'hC0, 8'hC0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h3E, 8'h60, 8'hC0, 8'hCE, 8'hC6, 8'h66, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC6, 8'hC6, 8'hC6, 8'hFE, 8'hC6, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h3C, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h1E, 8'h06, 8'h06, 8'h06, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC6, 8'hCC, 8'hD8, 8'hF0, 8'hD8, 8'hCC, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC6, 8'hEE, 8'hFE, 8'hFE, 8'hD6, 8'hC6, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC6, 8'hE6, 8'hF6, 8'hFE, 8'hDE, 8'hCE, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFC, 8'hC6, 8'hC6, 8'hFC, 8'hC0, 8'hC0, 8'hC0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h7C, 8'hC6, 8'hC6, 8'hC6, 8'hDE, 8'hCC, 8'h7A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFC, 8'hC6, 8'hC6, 8'hFC, 8'hD8, 8'hCC, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h78, 8'hCC, 8'hC0, 8'h7C, 8'h06, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h7E, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'hC6, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC6, 8'hC6, 8'hC6, 8'hEE, 8'h7C, 8'h38, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC6, 8'hC6, 8'hD6, 8'hFE, 8'hFE, 8'hEE, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hC6, 8'hEE, 8'h7C, 8'h38, 8'h7C, 8'hEE, 8'hC6, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h66, 8'h66, 8'h66, 8'h3C, 8'h18, 8'h18, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFE, 8'h0E, 8'h1C, 8'h38, 8'h70, 8'hE0, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h7E, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h18, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h6C, 8'h6C, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h7E, 8'h7E, 8'h00, 8'h7E, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h18, 8'h3C, 8'h3C, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h18, 8'h34, 8'h3C, 8'h18, 8'h08, 8'h10, 8'h00,
			8'h00, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h18, 8'h18, 8'h18, 8'h18, 8'h18, 8'h00, 8'h18, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h7C, 8'hC6, 8'h06, 8'h1C, 8'h30, 8'h00, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h92, 8'h54, 8'h38, 8'hFE, 8'h38, 8'h54, 8'h92, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h24, 8'h1A, 8'h65, 8'h90, 8'hDB, 8'h27, 8'h3F, 8'h1F, 8'h18, 8'h65, 8'h1A, 8'h6F, 8'h24, 8'h7B, 8'h3F, 8'h1F,
			8'h82, 8'h69, 8'h8A, 8'h25, 8'h5A, 8'hBF, 8'hFF, 8'hC3, 8'h4C, 8'h96, 8'h75, 8'hDA, 8'hA7, 8'hDF, 8'hFF, 8'hC3,
			8'h10, 8'hA5, 8'h50, 8'h4D, 8'hA2, 8'h8B, 8'hFF, 8'hE3, 8'h4C, 8'h5A, 8'hAF, 8'hB2, 8'h5D, 8'hF7, 8'hFF, 8'hE3,
			8'h34, 8'h4A, 8'hA6, 8'h28, 8'h52, 8'hC4, 8'hFC, 8'hF8, 8'h48, 8'hB4, 8'h58, 8'hD7, 8'hAD, 8'hBF, 8'hFE, 8'hF8,
			8'h0B, 8'h17, 8'h2F, 8'h17, 8'h0F, 8'h07, 8'h08, 8'h17, 8'h1F, 8'h3F, 8'h3F, 8'h3F, 8'h1F, 8'h0F, 8'h1F, 8'h1F,
			8'hF8, 8'hFC, 8'hFC, 8'hFC, 8'hF8, 8'hE0, 8'h18, 8'hF8, 8'hF8, 8'hFC, 8'hFC, 8'hFC, 8'hF8, 8'hF0, 8'hF8, 8'hF8,
			8'h0B, 8'h17, 8'h0B, 8'h05, 8'h03, 8'h00, 8'h00, 8'h00, 8'h1F, 8'h1F, 8'h0F, 8'h0F, 8'h07, 8'h00, 8'h00, 8'h00,
			8'hF8, 8'hF8, 8'hF0, 8'hF0, 8'hE0, 8'h00, 8'h00, 8'h00, 8'hF8, 8'hF8, 8'hF0, 8'hF0, 8'hE0, 8'h00, 8'h00, 8'h00,
			8'h82, 8'h69, 8'h8A, 8'h25, 8'h5A, 8'hBF, 8'hFF, 8'hFF, 8'h4C, 8'h96, 8'h75, 8'hDA, 8'hA7, 8'hDF, 8'hFF, 8'hFF,
			8'h10, 8'hA5, 8'h50, 8'h4D, 8'hA2, 8'h8B, 8'hFF, 8'hFF, 8'h4C, 8'h5A, 8'hAF, 8'hB2, 8'h5D, 8'hF7, 8'hFF, 8'hFF,
			8'h2F, 8'h1F, 8'h2F, 8'h5F, 8'hAF, 8'h5E, 8'hBC, 8'h18, 8'h3F, 8'h3F, 8'h7F, 8'h7F, 8'hFF, 8'hFE, 8'hFC, 8'h98,
			8'hBF, 8'h3B, 8'h59, 8'h3B, 8'h5F, 8'hBF, 8'h7E, 8'h0C, 8'hBF, 8'h7F, 8'h7B, 8'h7B, 8'h7F, 8'hFF, 8'h7E, 8'h0C,
			8'hFB, 8'hF5, 8'hD9, 8'h9C, 8'hBA, 8'hFC, 8'h3F, 8'h19, 8'hFF, 8'hFD, 8'hFD, 8'hDE, 8'hBE, 8'hFE, 8'h3F, 8'h19,
			8'hF8, 8'hF4, 8'hDA, 8'hDC, 8'hFA, 8'hFD, 8'h7E, 8'h01, 8'hFC, 8'hFC, 8'hDE, 8'hDE, 8'hFF, 8'hFF, 8'h7F, 8'h03,
			8'h24, 8'hAB, 8'h44, 8'hDB, 8'hFF, 8'hBF, 8'h5F, 8'h3C, 8'h5A, 8'h54, 8'hBB, 8'h3D, 8'hFF, 8'hFF, 8'h7F, 8'h7E,
			8'h42, 8'hBE, 8'h5F, 8'hBF, 8'h7F, 8'hBF, 8'h5F, 8'h3C, 8'h7E, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h7E,
			8'h42, 8'h3E, 8'h5E, 8'h2E, 8'h1E, 8'h3C, 8'h1C, 8'h08, 8'h7E, 8'h7E, 8'h7E, 8'h7E, 8'h3E, 8'h3C, 8'h3C, 8'h18,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'hDC, 8'h8F, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'hF8, 8'hFF, 8'hFF,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h8C, 8'h07, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'hF8, 8'hFB, 8'hFF,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'hDC, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hF8, 8'hFF, 8'hFF,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'hEC, 8'h87, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'hF8, 8'hFF, 8'hFF,
			8'h81, 8'h67, 8'h1E, 8'h04, 8'hC0, 8'h73, 8'h3A, 8'h10, 8'h7E, 8'hFD, 8'hFF, 8'hFF, 8'h3F, 8'hEF, 8'hFF, 8'hFF,
			8'h81, 8'h66, 8'h1C, 8'h18, 8'hC0, 8'h73, 8'h3C, 8'h00, 8'hFF, 8'hF9, 8'hFF, 8'hFF, 8'hBF, 8'hDF, 8'hFF, 8'hFF,
			8'h81, 8'h67, 8'h3E, 8'h08, 8'hC0, 8'h73, 8'h3D, 8'h18, 8'h7F, 8'hFB, 8'hF7, 8'hFF, 8'h7F, 8'hDF, 8'hFF, 8'hFF,
			8'h81, 8'h47, 8'h3E, 8'h04, 8'h40, 8'hF3, 8'h3D, 8'h08, 8'h7E, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hF7, 8'hFF,
			8'h81, 8'h47, 8'h36, 8'h0C, 8'hC0, 8'h73, 8'h3A, 8'h00, 8'h00, 8'hC5, 8'hFF, 8'hFF, 8'hBF, 8'hEF, 8'hFF, 8'hFF,
			8'h81, 8'h66, 8'h3F, 8'h02, 8'hC0, 8'h72, 8'h1C, 8'h08, 8'h80, 8'hE3, 8'hFD, 8'hFF, 8'hBF, 8'hDF, 8'hFF, 8'hFF,
			8'h81, 8'h67, 8'h3F, 8'h04, 8'hC0, 8'h73, 8'h3C, 8'h38, 8'h01, 8'hE5, 8'hFB, 8'hFF, 8'h3F, 8'hDF, 8'hEF, 8'hFF,
			8'h81, 8'h66, 8'h3C, 8'h1C, 8'hC0, 8'h72, 8'h3C, 8'h0C, 8'h00, 8'hE3, 8'hF7, 8'hFF, 8'h7F, 8'hDF, 8'hEF, 8'hFF,
			8'h00, 8'h00, 8'h01, 8'h03, 8'h03, 8'h03, 8'h07, 8'h07, 8'h03, 8'h07, 8'h0F, 8'h0E, 8'h1E, 8'h1E, 8'h1C, 8'h1C,
			8'h07, 8'h0B, 8'h0F, 8'h1F, 8'h3F, 8'h3F, 8'h7F, 8'h7D, 8'h08, 8'h1C, 8'h38, 8'h70, 8'h60, 8'hE1, 8'hC2, 8'hC2,
			8'hFD, 8'hFE, 8'hFE, 8'h7F, 8'h79, 8'h33, 8'h07, 8'h06, 8'hC2, 8'h81, 8'h81, 8'h00, 8'h46, 8'h3F, 8'h1F, 8'h1E,
			8'h0F, 8'h0F, 8'h0F, 8'h07, 8'h07, 8'h07, 8'h03, 8'h01, 8'h3C, 8'h3C, 8'h3C, 8'h1C, 8'h1C, 8'h0E, 8'h07, 8'h03,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h03, 8'h00, 8'h00, 8'h00, 8'h01, 8'h03, 8'h03, 8'h07, 8'h06,
			8'h3B, 8'h4F, 8'hF3, 8'hFD, 8'hFD, 8'hFD, 8'hFE, 8'hFE, 8'hC4, 8'hF0, 8'h8C, 8'h02, 8'h02, 8'h02, 8'h01, 8'h01,
			8'hFF, 8'hFF, 8'hFC, 8'h73, 8'h8F, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h80, 8'h8F, 8'hFC, 8'h70, 8'h80, 8'h00, 8'h00,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hDF, 8'hEF, 8'h00, 8'h00, 8'h00, 8'h06, 8'h0C, 8'h18, 8'h38, 8'hDC,
			8'h07, 8'h07, 8'h03, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h0E, 8'h07, 8'h07, 8'h03, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h07, 8'h0F, 8'h3F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h0F, 8'h3F, 8'hFF, 8'hF8, 8'hE0, 8'h80, 8'h00, 8'h00,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h01, 8'h01,
			8'hFE, 8'hFE, 8'hFC, 8'hF8, 8'h70, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h00, 8'h80, 8'hF0, 8'h00, 8'h00, 8'h00,
			8'h00, 8'hC0, 8'hF0, 8'hF8, 8'hFC, 8'hFE, 8'hFE, 8'hFF, 8'h00, 8'hC0, 8'hF0, 8'h38, 8'h0C, 8'h07, 8'h03, 8'h01,
			8'hFE, 8'hE1, 8'hDE, 8'hBF, 8'hBF, 8'hFF, 8'hFF, 8'hFF, 8'h1F, 8'h3E, 8'h61, 8'h40, 8'h40, 8'h00, 8'h00, 8'h00,
			8'hFF, 8'h7F, 8'h7F, 8'h3F, 8'h1F, 8'h0F, 8'h07, 8'h00, 8'h80, 8'hC0, 8'hC0, 8'h60, 8'h30, 8'h3C, 8'h0F, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h78, 8'hFC, 8'hFC, 8'hFE, 8'h00, 8'h00, 8'h00, 8'h78, 8'h8C, 8'h06, 8'h06, 8'h03,
			8'hFE, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h03, 8'h03, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hF0, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h40, 8'h30, 8'h1F, 8'h0F, 8'h00,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'hFE, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h02, 8'h01, 8'h00,
			8'hFE, 8'hFC, 8'hFC, 8'hF8, 8'hF8, 8'hF0, 8'hC0, 8'h00, 8'h02, 8'h04, 8'h04, 8'h00, 8'h08, 8'h30, 8'hC0, 8'h00,
			8'hE0, 8'h78, 8'hFC, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'h98, 8'h04, 8'h04, 8'h02, 8'h01, 8'h01, 8'h01,
			8'hFF, 8'hFF, 8'hDE, 8'hDC, 8'hB0, 8'h70, 8'hF8, 8'hFC, 8'h00, 8'h20, 8'h61, 8'h62, 8'hCC, 8'hB0, 8'h18, 8'h0C,
			8'hFC, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hF8, 8'hF0, 8'h04, 8'h06, 8'h02, 8'h02, 8'h02, 8'h02, 8'h04, 8'h08,
			8'hE8, 8'hFE, 8'hFE, 8'hFE, 8'hFC, 8'hFC, 8'hF8, 8'hE0, 8'h14, 8'h02, 8'h02, 8'h02, 8'h04, 8'h04, 8'h18, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h06, 8'h1F, 8'h3F, 8'h31, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h1F, 8'h1F,
			8'h60, 8'h60, 8'h21, 8'h11, 8'h31, 8'h79, 8'h61, 8'hC0, 8'h3F, 8'h3F, 8'h1E, 8'h0E, 8'h0F, 8'h17, 8'h3F, 8'h7F,
			8'h80, 8'h80, 8'h80, 8'h00, 8'h47, 8'h3F, 8'h1F, 8'h1E, 8'h7F, 8'h7F, 8'hFF, 8'h7F, 8'h79, 8'h33, 8'h07, 8'h07,
			8'h3C, 8'h3C, 8'h3C, 8'h1C, 8'h1C, 8'h0E, 8'h07, 8'h03, 8'h0F, 8'h0F, 8'h0F, 8'h07, 8'h07, 8'h07, 8'h03, 8'h01,
			8'h00, 8'h00, 8'h39, 8'h7F, 8'h66, 8'hC2, 8'hC0, 8'hF8, 8'h00, 8'h00, 8'h08, 8'h3D, 8'h7B, 8'h7F, 8'hBF, 8'hC7,
			8'hFC, 8'hF2, 8'hC0, 8'h80, 8'h80, 8'h00, 8'h00, 8'h80, 8'h1B, 8'h7D, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'h00, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'h02, 8'h14, 8'h0C, 8'h0E, 8'h0E, 8'h07, 8'h13, 8'hC0, 8'hFD, 8'hEB, 8'hF7, 8'hF7, 8'hF3, 8'hF1, 8'hF0, 8'hC0,
			8'h00, 8'h00, 8'hC0, 8'hE0, 8'h20, 8'h57, 8'h1E, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h80, 8'hC0, 8'hA1, 8'hE7, 8'hEF,
			8'h08, 8'h08, 8'h18, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hF7, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'h00, 8'h00, 8'h04, 8'h04, 8'hF8, 8'h70, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h77, 8'h8F, 8'hFF, 8'hFF,
			8'h00, 8'h04, 8'h02, 8'h01, 8'h04, 8'h08, 8'hE0, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFC, 8'hF8, 8'hE0, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'h60, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'hE0, 8'hF0,
			8'h00, 8'h08, 8'h00, 8'h00, 8'h08, 8'h18, 8'h7C, 8'h3E, 8'hF0, 8'hF8, 8'hF8, 8'hF8, 8'hF0, 8'hE0, 8'hD8, 8'hFC,
			8'h26, 8'h03, 8'h01, 8'h01, 8'h00, 8'h02, 8'h24, 8'h10, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hD8, 8'hE0,
			8'h10, 8'h00, 8'h20, 8'hC0, 8'h00, 8'h00, 8'h00, 8'h00, 8'hE0, 8'hE0, 8'hC0, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hF7, 8'hF7, 8'h25, 8'h25, 8'h25, 8'h25, 8'h27, 8'h27,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h70, 8'h70, 8'h50, 8'h56, 8'h76, 8'h70, 8'h40, 8'h40,
			8'hF0, 8'h60, 8'h60, 8'h66, 8'h66, 8'h60, 8'h60, 8'hF0, 8'hF0, 8'h60, 8'h60, 8'h66, 8'h66, 8'h60, 8'h60, 8'hF0,
			8'hF8, 8'h50, 8'h50, 8'h56, 8'h56, 8'h50, 8'h50, 8'hF8, 8'hF8, 8'h50, 8'h50, 8'h56, 8'h56, 8'h50, 8'h50, 8'hF8,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h20, 8'h40, 8'h40, 8'h40, 8'h40, 8'h20, 8'h10, 8'h00, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h3F, 8'h00,
			8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h1F, 8'h1F, 8'h1F, 8'h1F, 8'h1F, 8'h1F, 8'h1F, 8'h1F,
			8'h1C, 8'h0E, 8'h0E, 8'h0E, 8'h0E, 8'h1C, 8'h18, 8'h00, 8'hF6, 8'hFB, 8'hFB, 8'hFB, 8'hFB, 8'hF6, 8'hF4, 8'h00,
			8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'hD8, 8'hD8, 8'hD8, 8'hD8, 8'hD8, 8'hD8, 8'hD8, 8'hD8,
			8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'hFF,
			8'hC0, 8'h80, 8'h9F, 8'h9F, 8'h9F, 8'h80, 8'hC0, 8'hFF, 8'hC0, 8'h9F, 8'hBF, 8'hBF, 8'hBF, 8'h9F, 8'hC0, 8'hFF,
			8'h03, 8'h01, 8'hF9, 8'hF9, 8'hF9, 8'h01, 8'h03, 8'hFF, 8'h03, 8'hF9, 8'hFD, 8'hFD, 8'hFD, 8'hF9, 8'h03, 8'hFF,
			8'h00, 8'h3E, 8'h7F, 8'h7F, 8'h41, 8'h00, 8'h41, 8'h3E, 8'h00, 8'h3E, 8'h41, 8'h3E, 8'h7F, 8'h7F, 8'h7F, 8'h3E,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81, 8'h81, 8'h42, 8'h24, 8'h18, 8'h18, 8'h24, 8'h42, 8'h81,
			8'h1C, 8'h3E, 8'h7F, 8'h7F, 8'h7F, 8'h7F, 8'h3E, 8'h00, 8'h1C, 8'h3A, 8'h7B, 8'h7F, 8'h7F, 8'h7F, 8'h3E, 8'h1C,
			8'h0C, 8'h1C, 8'h00, 8'h18, 8'h10, 8'h00, 8'h38, 8'h30, 8'h00, 8'h10, 8'h3C, 8'h3C, 8'h34, 8'h3C, 8'h08, 8'h00,
			8'h00, 8'h7C, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'h7C, 8'h38, 8'h38, 8'h7C, 8'hFE, 8'hFE, 8'hBE, 8'hBE, 8'h7C, 8'h38,
			8'h00, 8'h00, 8'h07, 8'h0F, 8'h0F, 8'h1F, 8'h1F, 8'h1F, 8'h00, 8'h00, 8'h07, 8'h0C, 8'h0E, 8'h1F, 8'h1F, 8'h1F,
			8'h00, 8'h00, 8'h00, 8'h80, 8'h80, 8'hC0, 8'hC0, 8'h80, 8'h00, 8'h00, 8'h00, 8'h80, 8'h80, 8'hC0, 8'hC0, 8'hC0,
			8'h0F, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h07, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h40, 8'hF8, 8'h40, 8'h10, 8'h18, 8'h02, 8'h1F, 8'h02, 8'h80, 8'h18, 8'h3C, 8'h34, 8'h3C, 8'h3C, 8'h18, 8'h01,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h60, 8'hF0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hE0, 8'hF0,
			8'h01, 8'h03, 8'h03, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00, 8'h03, 8'h03, 8'h03, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00,
			8'hF8, 8'hF8, 8'hF8, 8'hF8, 8'hF0, 8'hE0, 8'h00, 8'h00, 8'hF8, 8'hF8, 8'hF8, 8'h78, 8'h30, 8'hE0, 8'h00, 8'h00,
			8'h38, 8'h7C, 8'hFD, 8'hFD, 8'hFC, 8'hFC, 8'h7C, 8'h38, 8'h38, 8'h5C, 8'hBE, 8'hFE, 8'hFE, 8'hFE, 8'h7C, 8'h38,
			8'h00, 8'h18, 8'hC0, 8'hCA, 8'h5B, 8'h03, 8'h18, 8'h00, 8'h00, 8'h18, 8'h3C, 8'h2E, 8'h7C, 8'h3C, 8'h18, 8'h00,
			8'h1C, 8'h3E, 8'h3F, 8'h3F, 8'hBF, 8'hBF, 8'h3E, 8'h1C, 8'h1C, 8'h3E, 8'h7F, 8'h7F, 8'h7F, 8'h7D, 8'h3A, 8'h1C,
			8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h03, 8'h03, 8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h03, 8'h03, 8'h03,
			8'h00, 8'h00, 8'hE0, 8'hF0, 8'hF8, 8'hF8, 8'hF8, 8'hF8, 8'h00, 8'h00, 8'hE0, 8'hF0, 8'hF8, 8'hF8, 8'hE8, 8'hC8,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0F,
			8'h02, 8'h1F, 8'h02, 8'h18, 8'h08, 8'h40, 8'hF8, 8'h40, 8'h01, 8'h18, 8'h3C, 8'h3C, 8'h2C, 8'h3C, 8'h18, 8'h80,
			8'hF0, 8'h60, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hF0, 8'hE0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h1F, 8'h1F, 8'h1F, 8'h1F, 8'h0F, 8'h07, 8'h00, 8'h00, 8'h13, 8'h17, 8'h1F, 8'h1F, 8'h0F, 8'h07, 8'h00, 8'h00,
			8'h80, 8'hC0, 8'hC0, 8'h80, 8'h80, 8'h00, 8'h00, 8'h00, 8'hC0, 8'hC0, 8'hC0, 8'h80, 8'h80, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h1F, 8'h3F, 8'h7F, 8'h7F, 8'hFF, 8'hFF,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'h00, 8'h00, 8'h00, 8'h60, 8'h30, 8'h18, 8'h08, 8'h08, 8'h00, 8'hC0, 8'hF0, 8'h98, 8'hCC, 8'hE4, 8'hF6, 8'hF6,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hC3, 8'h81, 8'h81, 8'h00, 8'h00, 8'h81, 8'h81, 8'hC3,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h7F, 8'h3F, 8'h1F, 8'h07,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'hFE, 8'hFC, 8'hFC, 8'hF8, 8'hF0, 8'hC0,
			8'h00, 8'h00, 8'h00, 8'h0C, 8'h04, 8'h06, 8'h02, 8'h02, 8'h00, 8'h3C, 8'h7E, 8'h72, 8'hFB, 8'hF9, 8'hFD, 8'hFD,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h1F,
			8'h00, 8'h00, 8'h18, 8'h0C, 8'h04, 8'h04, 8'h00, 8'h00, 8'h00, 8'hFC, 8'hE6, 8'hF2, 8'hFA, 8'hFA, 8'hFE, 8'hFC,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7E, 8'h7E, 8'h3C,
			8'h00, 8'h00, 8'h00, 8'h30, 8'h18, 8'h0C, 8'h04, 8'h04, 8'h00, 8'hE0, 8'hF8, 8'hCC, 8'hE6, 8'hF2, 8'hFB, 8'hFB,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h7B, 8'h7B, 8'h12, 8'h12, 8'h12, 8'h12, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h60, 8'hE0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hC3, 8'h81, 8'h81, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h81, 8'h81, 8'hC3, 8'hFF,
			8'h3C, 8'h42, 8'h99, 8'hA1, 8'hA1, 8'h99, 8'h42, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hC3, 8'h81, 8'h80, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h3F, 8'h1F, 8'h0F,
			8'hFC, 8'hC6, 8'hC6, 8'hFC, 8'hD8, 8'hCC, 8'hC6, 8'h00, 8'hFC, 8'hC6, 8'hC6, 8'hFC, 8'hD8, 8'hCC, 8'hC6, 8'h00,
			8'h38, 8'h6C, 8'hC6, 8'hC6, 8'hFE, 8'hC6, 8'hC6, 8'h00, 8'h38, 8'h6C, 8'hC6, 8'hC6, 8'hFE, 8'hC6, 8'hC6, 8'h00,
			8'hC6, 8'hE6, 8'hF6, 8'hFE, 8'hDE, 8'hCE, 8'hC6, 8'h00, 8'hC6, 8'hE6, 8'hF6, 8'hFE, 8'hDE, 8'hCE, 8'hC6, 8'h00,
			8'hC6, 8'hCC, 8'hD8, 8'hF0, 8'hD8, 8'hCC, 8'hC6, 8'h00, 8'hC6, 8'hCC, 8'hD8, 8'hF0, 8'hD8, 8'hCC, 8'hC6, 8'h00,
			8'h00, 8'h00, 8'h7E, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7E, 8'h7E, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
			8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF,
			8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF
		};
	end
	
	wire chip_select_prg = (I_prg_addr >= 16'h8000);
	
	assign O_ciram_a10 = I_chr_addr[11];
	assign O_ciram_a11 = 1'b0;
	assign O_ciram_ce = 1'b1;
	assign O_irq = 1'b1;
	
	always @(posedge I_clock)
	begin
		if (I_prg_wren & chip_select_prg)
			prg_bits[14' (I_prg_addr)] <= I_prg_data;
		
		if (chip_select_prg)
			O_prg_data <= prg_bits[14' (I_prg_addr)];
		else
			O_prg_data <= 8'hff;
		
		if (I_chr_wren)
			chr_bits[13' (I_chr_addr)] <= I_chr_data;
		O_chr_data <= chr_bits[13' (I_chr_addr)];
	end
endmodule