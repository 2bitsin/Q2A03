
	if (t0 | (o0 & o2 & o3 & o5 & o7 & t1 & ~o1 & ~o4 & ~o6) | (o0 & o2 & o3 & o5 & o7 & t2 & ~o1 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t1 & ~o0 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t2 & ~o0 & ~o4 & ~o6) | (o1 & o3 & o5 & o6 & o7 & t1 & ~o0 & ~o2 & ~o4) | (o3 & o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2) | (o0 & o2 & o3 & o7 & t1 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o3 & o7 & t2 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o5 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o6) | (o0 & o3 & o5 & o7 & t1 & ~o1 & ~o2 & ~o4 & ~o6) | (o1 & o2 & o3 & o7 & t1 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o3 & o7 & t2 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o5 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o6) | (o3 & o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o7) | (o3 & o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o6) | (o3 & o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o5) | (o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3) | (o4 & o5 & o6 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3) | (o0 & o2 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o5 & o7 & t1 & ~o0 & ~o2 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & t1 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o5 & t2 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o6 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o6 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o3 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o5 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o3 & o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o6 & ~o7) | (o3 & o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o5 & ~o7) | (o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o5 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o4 & o6 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o2 & o5 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o3 & o4 & t1 & ~o0 & ~o1 & ~o2 & ~o5 & ~o6 & ~o7) | (o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o5 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o4 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6) | (o4 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7) | (o4 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7) | (o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		G_addr = curr_pc;
	
	if (t0 | (o0 & o2 & o3 & o5 & o7 & t1 & ~o1 & ~o4 & ~o6) | (o0 & o2 & o3 & o5 & o7 & t2 & ~o1 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t1 & ~o0 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t2 & ~o0 & ~o4 & ~o6) | (o1 & o3 & o5 & o6 & o7 & t1 & ~o0 & ~o2 & ~o4) | (o3 & o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2) | (o0 & o2 & o3 & o7 & t1 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o5 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o6) | (o0 & o2 & o5 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o6) | (o0 & o3 & o5 & o7 & t1 & ~o1 & ~o2 & ~o4 & ~o6) | (o1 & o2 & o3 & o7 & t1 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o5 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o6) | (o1 & o2 & o5 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o6) | (o3 & o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o7) | (o3 & o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o6) | (o3 & o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o5) | (o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3) | (o4 & o5 & o6 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3) | (o4 & o5 & o6 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3) | (o0 & o2 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o5 & o7 & t1 & ~o0 & ~o2 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & t1 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o5 & t2 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o6 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o6 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o5 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o2 & o5 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o3 & o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o6 & ~o7) | (o3 & o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o5 & ~o7) | (o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o5 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o5 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o4 & o6 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o4 & o6 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o2 & o5 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o5 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o3 & o4 & t1 & ~o0 & ~o1 & ~o2 & ~o5 & ~o6 & ~o7) | (o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o5 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o5 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o4 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o4 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6) | (o4 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7) | (o4 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7) | (o4 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7) | (o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		G_rdwr = 1;
	
	if (o4 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7)
		next_cycle = (~curr_p[N_bit] ? (curr_cycle + 1) : 0);
	
	if (t0 | (o0 & o2 & o3 & o5 & o7 & t1 & ~o1 & ~o4 & ~o6) | (o0 & o2 & o3 & o5 & o7 & t2 & ~o1 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t1 & ~o0 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t2 & ~o0 & ~o4 & ~o6) | (o0 & o2 & o3 & o7 & t1 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o3 & o7 & t2 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o5 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o6) | (o0 & o3 & o5 & o7 & t1 & ~o1 & ~o2 & ~o4 & ~o6) | (o1 & o2 & o3 & o7 & t1 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o3 & o7 & t2 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o5 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o6) | (o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3) | (o0 & o2 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o5 & o7 & t1 & ~o0 & ~o2 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & t1 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o5 & t2 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o6 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o3 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o5 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o2 & o5 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o5 & o6 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6) | (o4 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7) | (o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		{next_pch, next_pcl} = curr_pc + 1;
	
	if ((o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3) | (o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o4 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7))
		{next_adh, next_adl} = {8'h00, G_rd_data} + (curr_pc + 1) - {7'h00, G_rd_data[7], 8'h00};
	
	if ((o4 & o5 & o6 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3) | (o4 & o5 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o6 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o4 & o5 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o4 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7))
		G_addr = {curr_pch, curr_adl};
	
	if ((o4 & o5 & o6 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3) | (o4 & o5 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o6 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o4 & o5 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o4 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7))
		{next_pch, next_pcl} = curr_ad;
	
	if ((o4 & o5 & o6 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3) | (o4 & o5 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o6 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o4 & o5 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o7 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o4 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7))
		next_cycle = ((curr_adh != curr_pch) ? (curr_cycle + 1) : 0);
	
	if ((o0 & o2 & o3 & o5 & o7 & t2 & ~o1 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t2 & ~o0 & ~o4 & ~o6) | (o1 & o3 & o5 & o6 & o7 & t1 & ~o0 & ~o2 & ~o4) | (o3 & o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2) | (o0 & o2 & o3 & o7 & t2 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o5 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o6) | (o0 & o3 & o5 & o7 & t1 & ~o1 & ~o2 & ~o4 & ~o6) | (o1 & o2 & o3 & o7 & t2 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o5 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o6) | (o3 & o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o7) | (o3 & o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o6) | (o3 & o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o5) | (o4 & o5 & o6 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3) | (o0 & o2 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o5 & o7 & t1 & ~o0 & ~o2 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & t2 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o6 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o5 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o3 & o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o6 & ~o7) | (o3 & o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o5 & ~o7) | (o4 & o5 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7) | (o4 & o5 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6) | (o4 & o6 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5) | (o2 & o5 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o3 & o4 & t1 & ~o0 & ~o1 & ~o2 & ~o5 & ~o6 & ~o7) | (o4 & o5 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7) | (o4 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7) | (o4 & o7 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6) | (o5 & o6 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6) | (o4 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6 & ~o7) | (o5 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		next_cycle = 0;
	
	if (o3 & o4 & t1 & ~o0 & ~o1 & ~o2 & ~o5 & ~o6 & ~o7)
		next_p = curr_p & ~C_mask;
	
	if (t0 | (o0 & o2 & o3 & o5 & o7 & t1 & ~o1 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t1 & ~o0 & ~o4 & ~o6) | (o0 & o2 & o3 & o7 & t1 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o5 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o6) | (o1 & o2 & o3 & o7 & t1 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o5 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o6) | (o0 & o2 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o2 & o3 & o5 & t1 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o6 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o5 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o2 & o5 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		next_cycle = curr_cycle + 1;
	
	if ((o0 & o2 & o3 & o5 & o7 & t1 & ~o1 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t1 & ~o0 & ~o4 & ~o6) | (o0 & o2 & o3 & o7 & t1 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o5 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o6) | (o1 & o2 & o3 & o7 & t1 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o5 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o6) | (o0 & o2 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o2 & o3 & o5 & t1 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o6 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o7 & t1 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o5 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o2 & o5 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		next_adl = G_rd_data;
	
	if ((o5 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		G_addr = {8'h01, curr_s};
	
	if ((o0 & o2 & o3 & o7 & t2 & ~o1 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o3 & o7 & t2 & ~o0 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o2 & o3 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o5 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		G_rdwr = 0;
	
	if (o5 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7)
		G_wr_data = curr_pch;
	
	if ((o5 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7) | (o5 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		next_s = curr_s - 1;
	
	if (o5 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7)
		G_wr_data = curr_pcl;
	
	if ((o0 & o2 & o3 & o5 & o7 & t2 & ~o1 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t2 & ~o0 & ~o4 & ~o6) | (o0 & o2 & o3 & o7 & t2 & ~o1 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o3 & o7 & t2 & ~o0 & ~o4 & ~o5 & ~o6) | (o2 & o3 & o5 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o6) | (o2 & o3 & o5 & t2 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o3 & o6 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o2 & o3 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o5 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		next_adh = G_rd_data;
	
	if ((o2 & o3 & o6 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o7) | (o5 & t5 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6 & ~o7))
		{next_pch, next_pcl} = next_ad;
	
	if ((o0 & o2 & o5 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o6) | (o1 & o2 & o5 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o6) | (o0 & o2 & o7 & t1 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t1 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o2 & o5 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o2 & o5 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o7 & t1 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6))
		next_adh = 0;
	
	if ((o0 & o2 & o5 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o6) | (o1 & o2 & o5 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o6) | (o0 & o2 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6) | (o2 & o5 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o2 & o5 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7) | (o2 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6))
		G_addr = curr_ad;
	
	if ((o2 & o3 & o5 & t2 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o5 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7))
		next_p[Z_bit] = (G_rd_data & curr_a) == 0;
	
	if ((o2 & o3 & o5 & t2 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o5 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7))
		next_p[V_bit] = G_rd_data[6];
	
	if ((o2 & o3 & o5 & t2 & ~o0 & ~o1 & ~o4 & ~o6 & ~o7) | (o2 & o5 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6 & ~o7))
		next_p[N_bit] = G_rd_data[7];
	
	if (o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6 & ~o7)
		next_cycle = (curr_p[N_bit] ? (curr_cycle + 1) : 0);
	
	if (o3 & o4 & o5 & t1 & ~o0 & ~o1 & ~o2 & ~o6 & ~o7)
		next_p = curr_p | C_mask;
	
	if (o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o7)
		next_cycle = (~curr_p[V_bit] ? (curr_cycle + 1) : 0);
	
	if (o3 & o4 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o5 & ~o7)
		next_p = curr_p & ~I_mask;
	
	if ((o5 & o6 & t2 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7) | (o5 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7))
		next_s = curr_s + 1;
	
	if (o5 & o6 & t3 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7)
		next_pcl = G_rd_data;
	
	if (o5 & o6 & t4 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o7)
		next_pch = G_rd_data;
	
	if (o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o7)
		next_cycle = (curr_p[V_bit] ? (curr_cycle + 1) : 0);
	
	if (o3 & o4 & o5 & o6 & t1 & ~o0 & ~o1 & ~o2 & ~o7)
		next_p = curr_p | I_mask;
	
	if ((o2 & o3 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o5 & ~o6) | (o2 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6))
		G_wr_data = curr_y;
	
	if ((o0 & o2 & o3 & o7 & t2 & ~o1 & ~o4 & ~o5 & ~o6) | (o0 & o2 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o5 & ~o6))
		G_wr_data = curr_a;
	
	if ((o1 & o2 & o3 & o7 & t2 & ~o0 & ~o4 & ~o5 & ~o6) | (o1 & o2 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o5 & ~o6))
		G_wr_data = curr_x;
	
	if (o4 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5 & ~o6)
		next_cycle = (~curr_p[C_bit] ? (curr_cycle + 1) : 0);
	
	if ((o2 & o3 & o5 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o6) | (o2 & o5 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6))
		next_y = G_rd_data;
	
	if ((o0 & o2 & o3 & o5 & o7 & t2 & ~o1 & ~o4 & ~o6) | (o1 & o2 & o3 & o5 & o7 & t2 & ~o0 & ~o4 & ~o6) | (o0 & o2 & o5 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o6) | (o0 & o3 & o5 & o7 & t1 & ~o1 & ~o2 & ~o4 & ~o6) | (o1 & o2 & o5 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o6) | (o2 & o3 & o5 & o7 & t2 & ~o0 & ~o1 & ~o4 & ~o6) | (o1 & o5 & o7 & t1 & ~o0 & ~o2 & ~o3 & ~o4 & ~o6) | (o2 & o5 & o7 & t2 & ~o0 & ~o1 & ~o3 & ~o4 & ~o6) | (o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o4 & ~o6))
		{next_p[N_bit], next_p[Z_bit]} = {G_rd_data[7], G_rd_data == 0};
	
	if ((o1 & o2 & o3 & o5 & o7 & t2 & ~o0 & ~o4 & ~o6) | (o1 & o2 & o5 & o7 & t2 & ~o0 & ~o3 & ~o4 & ~o6) | (o1 & o5 & o7 & t1 & ~o0 & ~o2 & ~o3 & ~o4 & ~o6))
		next_x = G_rd_data;
	
	if ((o0 & o2 & o3 & o5 & o7 & t2 & ~o1 & ~o4 & ~o6) | (o0 & o2 & o5 & o7 & t2 & ~o1 & ~o3 & ~o4 & ~o6) | (o0 & o3 & o5 & o7 & t1 & ~o1 & ~o2 & ~o4 & ~o6))
		next_a = G_rd_data;
	
	if (o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o6)
		next_cycle = (curr_p[C_bit] ? (curr_cycle + 1) : 0);
	
	if (o3 & o4 & o5 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o6)
		next_p = curr_p & ~V_mask;
	
	if (o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3 & ~o5)
		next_cycle = (~curr_p[Z_bit] ? (curr_cycle + 1) : 0);
	
	if (o3 & o4 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o5)
		next_p = curr_p & ~D_mask;
	
	if (o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2 & ~o3)
		next_cycle = (curr_p[Z_bit] ? (curr_cycle + 1) : 0);
	
	if (o3 & o4 & o5 & o6 & o7 & t1 & ~o0 & ~o1 & ~o2)
		next_p = curr_p | D_mask;
	
	if (t0)
		next_ir = G_rd_data;
	