
module font8x16 (clock, addr, data);
	input wire clock;
	input wire[11:0] addr;
	output bit[7:0] data;
	always @(posedge clock)
	begin
		case(addr)
			12'h00000000 : data <= 8'b00000000 ;
			12'h00000001 : data <= 8'b00000000 ;
			12'h00000002 : data <= 8'b00000000 ;
			12'h00000003 : data <= 8'b00000000 ;
			12'h00000004 : data <= 8'b00000000 ;
			12'h00000005 : data <= 8'b00000000 ;
			12'h00000006 : data <= 8'b00000000 ;
			12'h00000007 : data <= 8'b00000000 ;
			12'h00000008 : data <= 8'b00000000 ;
			12'h00000009 : data <= 8'b00000000 ;
			12'h0000000A : data <= 8'b00000000 ;
			12'h0000000B : data <= 8'b00000000 ;
			12'h0000000C : data <= 8'b00000000 ;
			12'h0000000D : data <= 8'b00000000 ;
			12'h0000000E : data <= 8'b00000000 ;
			12'h0000000F : data <= 8'b00000000 ;
			12'h00000010 : data <= 8'b00000000 ;
			12'h00000011 : data <= 8'b00000000 ;
			12'h00000012 : data <= 8'b01111110 ;
			12'h00000013 : data <= 8'b10000001 ;
			12'h00000014 : data <= 8'b10100101 ;
			12'h00000015 : data <= 8'b10000001 ;
			12'h00000016 : data <= 8'b10000001 ;
			12'h00000017 : data <= 8'b10111101 ;
			12'h00000018 : data <= 8'b10011001 ;
			12'h00000019 : data <= 8'b10000001 ;
			12'h0000001A : data <= 8'b10000001 ;
			12'h0000001B : data <= 8'b01111110 ;
			12'h0000001C : data <= 8'b00000000 ;
			12'h0000001D : data <= 8'b00000000 ;
			12'h0000001E : data <= 8'b00000000 ;
			12'h0000001F : data <= 8'b00000000 ;
			12'h00000020 : data <= 8'b00000000 ;
			12'h00000021 : data <= 8'b00000000 ;
			12'h00000022 : data <= 8'b01111110 ;
			12'h00000023 : data <= 8'b11111111 ;
			12'h00000024 : data <= 8'b11011011 ;
			12'h00000025 : data <= 8'b11111111 ;
			12'h00000026 : data <= 8'b11111111 ;
			12'h00000027 : data <= 8'b11000011 ;
			12'h00000028 : data <= 8'b11100111 ;
			12'h00000029 : data <= 8'b11111111 ;
			12'h0000002A : data <= 8'b11111111 ;
			12'h0000002B : data <= 8'b01111110 ;
			12'h0000002C : data <= 8'b00000000 ;
			12'h0000002D : data <= 8'b00000000 ;
			12'h0000002E : data <= 8'b00000000 ;
			12'h0000002F : data <= 8'b00000000 ;
			12'h00000030 : data <= 8'b00000000 ;
			12'h00000031 : data <= 8'b00000000 ;
			12'h00000032 : data <= 8'b00000000 ;
			12'h00000033 : data <= 8'b00000000 ;
			12'h00000034 : data <= 8'b01101100 ;
			12'h00000035 : data <= 8'b11111110 ;
			12'h00000036 : data <= 8'b11111110 ;
			12'h00000037 : data <= 8'b11111110 ;
			12'h00000038 : data <= 8'b11111110 ;
			12'h00000039 : data <= 8'b01111100 ;
			12'h0000003A : data <= 8'b00111000 ;
			12'h0000003B : data <= 8'b00010000 ;
			12'h0000003C : data <= 8'b00000000 ;
			12'h0000003D : data <= 8'b00000000 ;
			12'h0000003E : data <= 8'b00000000 ;
			12'h0000003F : data <= 8'b00000000 ;
			12'h00000040 : data <= 8'b00000000 ;
			12'h00000041 : data <= 8'b00000000 ;
			12'h00000042 : data <= 8'b00000000 ;
			12'h00000043 : data <= 8'b00000000 ;
			12'h00000044 : data <= 8'b00010000 ;
			12'h00000045 : data <= 8'b00111000 ;
			12'h00000046 : data <= 8'b01111100 ;
			12'h00000047 : data <= 8'b11111110 ;
			12'h00000048 : data <= 8'b01111100 ;
			12'h00000049 : data <= 8'b00111000 ;
			12'h0000004A : data <= 8'b00010000 ;
			12'h0000004B : data <= 8'b00000000 ;
			12'h0000004C : data <= 8'b00000000 ;
			12'h0000004D : data <= 8'b00000000 ;
			12'h0000004E : data <= 8'b00000000 ;
			12'h0000004F : data <= 8'b00000000 ;
			12'h00000050 : data <= 8'b00000000 ;
			12'h00000051 : data <= 8'b00000000 ;
			12'h00000052 : data <= 8'b00000000 ;
			12'h00000053 : data <= 8'b00011000 ;
			12'h00000054 : data <= 8'b00111100 ;
			12'h00000055 : data <= 8'b00111100 ;
			12'h00000056 : data <= 8'b11100111 ;
			12'h00000057 : data <= 8'b11100111 ;
			12'h00000058 : data <= 8'b11100111 ;
			12'h00000059 : data <= 8'b00011000 ;
			12'h0000005A : data <= 8'b00011000 ;
			12'h0000005B : data <= 8'b00111100 ;
			12'h0000005C : data <= 8'b00000000 ;
			12'h0000005D : data <= 8'b00000000 ;
			12'h0000005E : data <= 8'b00000000 ;
			12'h0000005F : data <= 8'b00000000 ;
			12'h00000060 : data <= 8'b00000000 ;
			12'h00000061 : data <= 8'b00000000 ;
			12'h00000062 : data <= 8'b00000000 ;
			12'h00000063 : data <= 8'b00011000 ;
			12'h00000064 : data <= 8'b00111100 ;
			12'h00000065 : data <= 8'b01111110 ;
			12'h00000066 : data <= 8'b11111111 ;
			12'h00000067 : data <= 8'b11111111 ;
			12'h00000068 : data <= 8'b01111110 ;
			12'h00000069 : data <= 8'b00011000 ;
			12'h0000006A : data <= 8'b00011000 ;
			12'h0000006B : data <= 8'b00111100 ;
			12'h0000006C : data <= 8'b00000000 ;
			12'h0000006D : data <= 8'b00000000 ;
			12'h0000006E : data <= 8'b00000000 ;
			12'h0000006F : data <= 8'b00000000 ;
			12'h00000070 : data <= 8'b00000000 ;
			12'h00000071 : data <= 8'b00000000 ;
			12'h00000072 : data <= 8'b00000000 ;
			12'h00000073 : data <= 8'b00000000 ;
			12'h00000074 : data <= 8'b00000000 ;
			12'h00000075 : data <= 8'b00000000 ;
			12'h00000076 : data <= 8'b00011000 ;
			12'h00000077 : data <= 8'b00111100 ;
			12'h00000078 : data <= 8'b00111100 ;
			12'h00000079 : data <= 8'b00011000 ;
			12'h0000007A : data <= 8'b00000000 ;
			12'h0000007B : data <= 8'b00000000 ;
			12'h0000007C : data <= 8'b00000000 ;
			12'h0000007D : data <= 8'b00000000 ;
			12'h0000007E : data <= 8'b00000000 ;
			12'h0000007F : data <= 8'b00000000 ;
			12'h00000080 : data <= 8'b11111111 ;
			12'h00000081 : data <= 8'b11111111 ;
			12'h00000082 : data <= 8'b11111111 ;
			12'h00000083 : data <= 8'b11111111 ;
			12'h00000084 : data <= 8'b11111111 ;
			12'h00000085 : data <= 8'b11111111 ;
			12'h00000086 : data <= 8'b11100111 ;
			12'h00000087 : data <= 8'b11000011 ;
			12'h00000088 : data <= 8'b11000011 ;
			12'h00000089 : data <= 8'b11100111 ;
			12'h0000008A : data <= 8'b11111111 ;
			12'h0000008B : data <= 8'b11111111 ;
			12'h0000008C : data <= 8'b11111111 ;
			12'h0000008D : data <= 8'b11111111 ;
			12'h0000008E : data <= 8'b11111111 ;
			12'h0000008F : data <= 8'b11111111 ;
			12'h00000090 : data <= 8'b00000000 ;
			12'h00000091 : data <= 8'b00000000 ;
			12'h00000092 : data <= 8'b00000000 ;
			12'h00000093 : data <= 8'b00000000 ;
			12'h00000094 : data <= 8'b00000000 ;
			12'h00000095 : data <= 8'b00111100 ;
			12'h00000096 : data <= 8'b01100110 ;
			12'h00000097 : data <= 8'b01000010 ;
			12'h00000098 : data <= 8'b01000010 ;
			12'h00000099 : data <= 8'b01100110 ;
			12'h0000009A : data <= 8'b00111100 ;
			12'h0000009B : data <= 8'b00000000 ;
			12'h0000009C : data <= 8'b00000000 ;
			12'h0000009D : data <= 8'b00000000 ;
			12'h0000009E : data <= 8'b00000000 ;
			12'h0000009F : data <= 8'b00000000 ;
			12'h000000A0 : data <= 8'b11111111 ;
			12'h000000A1 : data <= 8'b11111111 ;
			12'h000000A2 : data <= 8'b11111111 ;
			12'h000000A3 : data <= 8'b11111111 ;
			12'h000000A4 : data <= 8'b11111111 ;
			12'h000000A5 : data <= 8'b11000011 ;
			12'h000000A6 : data <= 8'b10011001 ;
			12'h000000A7 : data <= 8'b10111101 ;
			12'h000000A8 : data <= 8'b10111101 ;
			12'h000000A9 : data <= 8'b10011001 ;
			12'h000000AA : data <= 8'b11000011 ;
			12'h000000AB : data <= 8'b11111111 ;
			12'h000000AC : data <= 8'b11111111 ;
			12'h000000AD : data <= 8'b11111111 ;
			12'h000000AE : data <= 8'b11111111 ;
			12'h000000AF : data <= 8'b11111111 ;
			12'h000000B0 : data <= 8'b00000000 ;
			12'h000000B1 : data <= 8'b00000000 ;
			12'h000000B2 : data <= 8'b00011110 ;
			12'h000000B3 : data <= 8'b00001110 ;
			12'h000000B4 : data <= 8'b00011010 ;
			12'h000000B5 : data <= 8'b00110010 ;
			12'h000000B6 : data <= 8'b01111000 ;
			12'h000000B7 : data <= 8'b11001100 ;
			12'h000000B8 : data <= 8'b11001100 ;
			12'h000000B9 : data <= 8'b11001100 ;
			12'h000000BA : data <= 8'b11001100 ;
			12'h000000BB : data <= 8'b01111000 ;
			12'h000000BC : data <= 8'b00000000 ;
			12'h000000BD : data <= 8'b00000000 ;
			12'h000000BE : data <= 8'b00000000 ;
			12'h000000BF : data <= 8'b00000000 ;
			12'h000000C0 : data <= 8'b00000000 ;
			12'h000000C1 : data <= 8'b00000000 ;
			12'h000000C2 : data <= 8'b00111100 ;
			12'h000000C3 : data <= 8'b01100110 ;
			12'h000000C4 : data <= 8'b01100110 ;
			12'h000000C5 : data <= 8'b01100110 ;
			12'h000000C6 : data <= 8'b01100110 ;
			12'h000000C7 : data <= 8'b00111100 ;
			12'h000000C8 : data <= 8'b00011000 ;
			12'h000000C9 : data <= 8'b01111110 ;
			12'h000000CA : data <= 8'b00011000 ;
			12'h000000CB : data <= 8'b00011000 ;
			12'h000000CC : data <= 8'b00000000 ;
			12'h000000CD : data <= 8'b00000000 ;
			12'h000000CE : data <= 8'b00000000 ;
			12'h000000CF : data <= 8'b00000000 ;
			12'h000000D0 : data <= 8'b00000000 ;
			12'h000000D1 : data <= 8'b00000000 ;
			12'h000000D2 : data <= 8'b00111111 ;
			12'h000000D3 : data <= 8'b00110011 ;
			12'h000000D4 : data <= 8'b00111111 ;
			12'h000000D5 : data <= 8'b00110000 ;
			12'h000000D6 : data <= 8'b00110000 ;
			12'h000000D7 : data <= 8'b00110000 ;
			12'h000000D8 : data <= 8'b00110000 ;
			12'h000000D9 : data <= 8'b01110000 ;
			12'h000000DA : data <= 8'b11110000 ;
			12'h000000DB : data <= 8'b11100000 ;
			12'h000000DC : data <= 8'b00000000 ;
			12'h000000DD : data <= 8'b00000000 ;
			12'h000000DE : data <= 8'b00000000 ;
			12'h000000DF : data <= 8'b00000000 ;
			12'h000000E0 : data <= 8'b00000000 ;
			12'h000000E1 : data <= 8'b00000000 ;
			12'h000000E2 : data <= 8'b01111111 ;
			12'h000000E3 : data <= 8'b01100011 ;
			12'h000000E4 : data <= 8'b01111111 ;
			12'h000000E5 : data <= 8'b01100011 ;
			12'h000000E6 : data <= 8'b01100011 ;
			12'h000000E7 : data <= 8'b01100011 ;
			12'h000000E8 : data <= 8'b01100011 ;
			12'h000000E9 : data <= 8'b01100111 ;
			12'h000000EA : data <= 8'b11100111 ;
			12'h000000EB : data <= 8'b11100110 ;
			12'h000000EC : data <= 8'b11000000 ;
			12'h000000ED : data <= 8'b00000000 ;
			12'h000000EE : data <= 8'b00000000 ;
			12'h000000EF : data <= 8'b00000000 ;
			12'h000000F0 : data <= 8'b00000000 ;
			12'h000000F1 : data <= 8'b00000000 ;
			12'h000000F2 : data <= 8'b00000000 ;
			12'h000000F3 : data <= 8'b00011000 ;
			12'h000000F4 : data <= 8'b00011000 ;
			12'h000000F5 : data <= 8'b11011011 ;
			12'h000000F6 : data <= 8'b00111100 ;
			12'h000000F7 : data <= 8'b11100111 ;
			12'h000000F8 : data <= 8'b00111100 ;
			12'h000000F9 : data <= 8'b11011011 ;
			12'h000000FA : data <= 8'b00011000 ;
			12'h000000FB : data <= 8'b00011000 ;
			12'h000000FC : data <= 8'b00000000 ;
			12'h000000FD : data <= 8'b00000000 ;
			12'h000000FE : data <= 8'b00000000 ;
			12'h000000FF : data <= 8'b00000000 ;
			12'h00000100 : data <= 8'b00000000 ;
			12'h00000101 : data <= 8'b10000000 ;
			12'h00000102 : data <= 8'b11000000 ;
			12'h00000103 : data <= 8'b11100000 ;
			12'h00000104 : data <= 8'b11110000 ;
			12'h00000105 : data <= 8'b11111000 ;
			12'h00000106 : data <= 8'b11111110 ;
			12'h00000107 : data <= 8'b11111000 ;
			12'h00000108 : data <= 8'b11110000 ;
			12'h00000109 : data <= 8'b11100000 ;
			12'h0000010A : data <= 8'b11000000 ;
			12'h0000010B : data <= 8'b10000000 ;
			12'h0000010C : data <= 8'b00000000 ;
			12'h0000010D : data <= 8'b00000000 ;
			12'h0000010E : data <= 8'b00000000 ;
			12'h0000010F : data <= 8'b00000000 ;
			12'h00000110 : data <= 8'b00000000 ;
			12'h00000111 : data <= 8'b00000010 ;
			12'h00000112 : data <= 8'b00000110 ;
			12'h00000113 : data <= 8'b00001110 ;
			12'h00000114 : data <= 8'b00011110 ;
			12'h00000115 : data <= 8'b00111110 ;
			12'h00000116 : data <= 8'b11111110 ;
			12'h00000117 : data <= 8'b00111110 ;
			12'h00000118 : data <= 8'b00011110 ;
			12'h00000119 : data <= 8'b00001110 ;
			12'h0000011A : data <= 8'b00000110 ;
			12'h0000011B : data <= 8'b00000010 ;
			12'h0000011C : data <= 8'b00000000 ;
			12'h0000011D : data <= 8'b00000000 ;
			12'h0000011E : data <= 8'b00000000 ;
			12'h0000011F : data <= 8'b00000000 ;
			12'h00000120 : data <= 8'b00000000 ;
			12'h00000121 : data <= 8'b00000000 ;
			12'h00000122 : data <= 8'b00011000 ;
			12'h00000123 : data <= 8'b00111100 ;
			12'h00000124 : data <= 8'b01111110 ;
			12'h00000125 : data <= 8'b00011000 ;
			12'h00000126 : data <= 8'b00011000 ;
			12'h00000127 : data <= 8'b00011000 ;
			12'h00000128 : data <= 8'b01111110 ;
			12'h00000129 : data <= 8'b00111100 ;
			12'h0000012A : data <= 8'b00011000 ;
			12'h0000012B : data <= 8'b00000000 ;
			12'h0000012C : data <= 8'b00000000 ;
			12'h0000012D : data <= 8'b00000000 ;
			12'h0000012E : data <= 8'b00000000 ;
			12'h0000012F : data <= 8'b00000000 ;
			12'h00000130 : data <= 8'b00000000 ;
			12'h00000131 : data <= 8'b00000000 ;
			12'h00000132 : data <= 8'b01100110 ;
			12'h00000133 : data <= 8'b01100110 ;
			12'h00000134 : data <= 8'b01100110 ;
			12'h00000135 : data <= 8'b01100110 ;
			12'h00000136 : data <= 8'b01100110 ;
			12'h00000137 : data <= 8'b01100110 ;
			12'h00000138 : data <= 8'b01100110 ;
			12'h00000139 : data <= 8'b00000000 ;
			12'h0000013A : data <= 8'b01100110 ;
			12'h0000013B : data <= 8'b01100110 ;
			12'h0000013C : data <= 8'b00000000 ;
			12'h0000013D : data <= 8'b00000000 ;
			12'h0000013E : data <= 8'b00000000 ;
			12'h0000013F : data <= 8'b00000000 ;
			12'h00000140 : data <= 8'b00000000 ;
			12'h00000141 : data <= 8'b00000000 ;
			12'h00000142 : data <= 8'b01111111 ;
			12'h00000143 : data <= 8'b11011011 ;
			12'h00000144 : data <= 8'b11011011 ;
			12'h00000145 : data <= 8'b11011011 ;
			12'h00000146 : data <= 8'b01111011 ;
			12'h00000147 : data <= 8'b00011011 ;
			12'h00000148 : data <= 8'b00011011 ;
			12'h00000149 : data <= 8'b00011011 ;
			12'h0000014A : data <= 8'b00011011 ;
			12'h0000014B : data <= 8'b00011011 ;
			12'h0000014C : data <= 8'b00000000 ;
			12'h0000014D : data <= 8'b00000000 ;
			12'h0000014E : data <= 8'b00000000 ;
			12'h0000014F : data <= 8'b00000000 ;
			12'h00000150 : data <= 8'b00000000 ;
			12'h00000151 : data <= 8'b01111100 ;
			12'h00000152 : data <= 8'b11000110 ;
			12'h00000153 : data <= 8'b01100000 ;
			12'h00000154 : data <= 8'b00111000 ;
			12'h00000155 : data <= 8'b01101100 ;
			12'h00000156 : data <= 8'b11000110 ;
			12'h00000157 : data <= 8'b11000110 ;
			12'h00000158 : data <= 8'b01101100 ;
			12'h00000159 : data <= 8'b00111000 ;
			12'h0000015A : data <= 8'b00001100 ;
			12'h0000015B : data <= 8'b11000110 ;
			12'h0000015C : data <= 8'b01111100 ;
			12'h0000015D : data <= 8'b00000000 ;
			12'h0000015E : data <= 8'b00000000 ;
			12'h0000015F : data <= 8'b00000000 ;
			12'h00000160 : data <= 8'b00000000 ;
			12'h00000161 : data <= 8'b00000000 ;
			12'h00000162 : data <= 8'b00000000 ;
			12'h00000163 : data <= 8'b00000000 ;
			12'h00000164 : data <= 8'b00000000 ;
			12'h00000165 : data <= 8'b00000000 ;
			12'h00000166 : data <= 8'b00000000 ;
			12'h00000167 : data <= 8'b00000000 ;
			12'h00000168 : data <= 8'b11111110 ;
			12'h00000169 : data <= 8'b11111110 ;
			12'h0000016A : data <= 8'b11111110 ;
			12'h0000016B : data <= 8'b11111110 ;
			12'h0000016C : data <= 8'b00000000 ;
			12'h0000016D : data <= 8'b00000000 ;
			12'h0000016E : data <= 8'b00000000 ;
			12'h0000016F : data <= 8'b00000000 ;
			12'h00000170 : data <= 8'b00000000 ;
			12'h00000171 : data <= 8'b00000000 ;
			12'h00000172 : data <= 8'b00011000 ;
			12'h00000173 : data <= 8'b00111100 ;
			12'h00000174 : data <= 8'b01111110 ;
			12'h00000175 : data <= 8'b00011000 ;
			12'h00000176 : data <= 8'b00011000 ;
			12'h00000177 : data <= 8'b00011000 ;
			12'h00000178 : data <= 8'b01111110 ;
			12'h00000179 : data <= 8'b00111100 ;
			12'h0000017A : data <= 8'b00011000 ;
			12'h0000017B : data <= 8'b01111110 ;
			12'h0000017C : data <= 8'b00000000 ;
			12'h0000017D : data <= 8'b00000000 ;
			12'h0000017E : data <= 8'b00000000 ;
			12'h0000017F : data <= 8'b00000000 ;
			12'h00000180 : data <= 8'b00000000 ;
			12'h00000181 : data <= 8'b00000000 ;
			12'h00000182 : data <= 8'b00011000 ;
			12'h00000183 : data <= 8'b00111100 ;
			12'h00000184 : data <= 8'b01111110 ;
			12'h00000185 : data <= 8'b00011000 ;
			12'h00000186 : data <= 8'b00011000 ;
			12'h00000187 : data <= 8'b00011000 ;
			12'h00000188 : data <= 8'b00011000 ;
			12'h00000189 : data <= 8'b00011000 ;
			12'h0000018A : data <= 8'b00011000 ;
			12'h0000018B : data <= 8'b00011000 ;
			12'h0000018C : data <= 8'b00000000 ;
			12'h0000018D : data <= 8'b00000000 ;
			12'h0000018E : data <= 8'b00000000 ;
			12'h0000018F : data <= 8'b00000000 ;
			12'h00000190 : data <= 8'b00000000 ;
			12'h00000191 : data <= 8'b00000000 ;
			12'h00000192 : data <= 8'b00011000 ;
			12'h00000193 : data <= 8'b00011000 ;
			12'h00000194 : data <= 8'b00011000 ;
			12'h00000195 : data <= 8'b00011000 ;
			12'h00000196 : data <= 8'b00011000 ;
			12'h00000197 : data <= 8'b00011000 ;
			12'h00000198 : data <= 8'b00011000 ;
			12'h00000199 : data <= 8'b01111110 ;
			12'h0000019A : data <= 8'b00111100 ;
			12'h0000019B : data <= 8'b00011000 ;
			12'h0000019C : data <= 8'b00000000 ;
			12'h0000019D : data <= 8'b00000000 ;
			12'h0000019E : data <= 8'b00000000 ;
			12'h0000019F : data <= 8'b00000000 ;
			12'h000001A0 : data <= 8'b00000000 ;
			12'h000001A1 : data <= 8'b00000000 ;
			12'h000001A2 : data <= 8'b00000000 ;
			12'h000001A3 : data <= 8'b00000000 ;
			12'h000001A4 : data <= 8'b00000000 ;
			12'h000001A5 : data <= 8'b00011000 ;
			12'h000001A6 : data <= 8'b00001100 ;
			12'h000001A7 : data <= 8'b11111110 ;
			12'h000001A8 : data <= 8'b00001100 ;
			12'h000001A9 : data <= 8'b00011000 ;
			12'h000001AA : data <= 8'b00000000 ;
			12'h000001AB : data <= 8'b00000000 ;
			12'h000001AC : data <= 8'b00000000 ;
			12'h000001AD : data <= 8'b00000000 ;
			12'h000001AE : data <= 8'b00000000 ;
			12'h000001AF : data <= 8'b00000000 ;
			12'h000001B0 : data <= 8'b00000000 ;
			12'h000001B1 : data <= 8'b00000000 ;
			12'h000001B2 : data <= 8'b00000000 ;
			12'h000001B3 : data <= 8'b00000000 ;
			12'h000001B4 : data <= 8'b00000000 ;
			12'h000001B5 : data <= 8'b00110000 ;
			12'h000001B6 : data <= 8'b01100000 ;
			12'h000001B7 : data <= 8'b11111110 ;
			12'h000001B8 : data <= 8'b01100000 ;
			12'h000001B9 : data <= 8'b00110000 ;
			12'h000001BA : data <= 8'b00000000 ;
			12'h000001BB : data <= 8'b00000000 ;
			12'h000001BC : data <= 8'b00000000 ;
			12'h000001BD : data <= 8'b00000000 ;
			12'h000001BE : data <= 8'b00000000 ;
			12'h000001BF : data <= 8'b00000000 ;
			12'h000001C0 : data <= 8'b00000000 ;
			12'h000001C1 : data <= 8'b00000000 ;
			12'h000001C2 : data <= 8'b00000000 ;
			12'h000001C3 : data <= 8'b00000000 ;
			12'h000001C4 : data <= 8'b00000000 ;
			12'h000001C5 : data <= 8'b00000000 ;
			12'h000001C6 : data <= 8'b11000000 ;
			12'h000001C7 : data <= 8'b11000000 ;
			12'h000001C8 : data <= 8'b11000000 ;
			12'h000001C9 : data <= 8'b11111110 ;
			12'h000001CA : data <= 8'b00000000 ;
			12'h000001CB : data <= 8'b00000000 ;
			12'h000001CC : data <= 8'b00000000 ;
			12'h000001CD : data <= 8'b00000000 ;
			12'h000001CE : data <= 8'b00000000 ;
			12'h000001CF : data <= 8'b00000000 ;
			12'h000001D0 : data <= 8'b00000000 ;
			12'h000001D1 : data <= 8'b00000000 ;
			12'h000001D2 : data <= 8'b00000000 ;
			12'h000001D3 : data <= 8'b00000000 ;
			12'h000001D4 : data <= 8'b00000000 ;
			12'h000001D5 : data <= 8'b00101000 ;
			12'h000001D6 : data <= 8'b01101100 ;
			12'h000001D7 : data <= 8'b11111110 ;
			12'h000001D8 : data <= 8'b01101100 ;
			12'h000001D9 : data <= 8'b00101000 ;
			12'h000001DA : data <= 8'b00000000 ;
			12'h000001DB : data <= 8'b00000000 ;
			12'h000001DC : data <= 8'b00000000 ;
			12'h000001DD : data <= 8'b00000000 ;
			12'h000001DE : data <= 8'b00000000 ;
			12'h000001DF : data <= 8'b00000000 ;
			12'h000001E0 : data <= 8'b00000000 ;
			12'h000001E1 : data <= 8'b00000000 ;
			12'h000001E2 : data <= 8'b00000000 ;
			12'h000001E3 : data <= 8'b00000000 ;
			12'h000001E4 : data <= 8'b00010000 ;
			12'h000001E5 : data <= 8'b00111000 ;
			12'h000001E6 : data <= 8'b00111000 ;
			12'h000001E7 : data <= 8'b01111100 ;
			12'h000001E8 : data <= 8'b01111100 ;
			12'h000001E9 : data <= 8'b11111110 ;
			12'h000001EA : data <= 8'b11111110 ;
			12'h000001EB : data <= 8'b00000000 ;
			12'h000001EC : data <= 8'b00000000 ;
			12'h000001ED : data <= 8'b00000000 ;
			12'h000001EE : data <= 8'b00000000 ;
			12'h000001EF : data <= 8'b00000000 ;
			12'h000001F0 : data <= 8'b00000000 ;
			12'h000001F1 : data <= 8'b00000000 ;
			12'h000001F2 : data <= 8'b00000000 ;
			12'h000001F3 : data <= 8'b00000000 ;
			12'h000001F4 : data <= 8'b11111110 ;
			12'h000001F5 : data <= 8'b11111110 ;
			12'h000001F6 : data <= 8'b01111100 ;
			12'h000001F7 : data <= 8'b01111100 ;
			12'h000001F8 : data <= 8'b00111000 ;
			12'h000001F9 : data <= 8'b00111000 ;
			12'h000001FA : data <= 8'b00010000 ;
			12'h000001FB : data <= 8'b00000000 ;
			12'h000001FC : data <= 8'b00000000 ;
			12'h000001FD : data <= 8'b00000000 ;
			12'h000001FE : data <= 8'b00000000 ;
			12'h000001FF : data <= 8'b00000000 ;
			12'h00000200 : data <= 8'b00000000 ;
			12'h00000201 : data <= 8'b00000000 ;
			12'h00000202 : data <= 8'b00000000 ;
			12'h00000203 : data <= 8'b00000000 ;
			12'h00000204 : data <= 8'b00000000 ;
			12'h00000205 : data <= 8'b00000000 ;
			12'h00000206 : data <= 8'b00000000 ;
			12'h00000207 : data <= 8'b00000000 ;
			12'h00000208 : data <= 8'b00000000 ;
			12'h00000209 : data <= 8'b00000000 ;
			12'h0000020A : data <= 8'b00000000 ;
			12'h0000020B : data <= 8'b00000000 ;
			12'h0000020C : data <= 8'b00000000 ;
			12'h0000020D : data <= 8'b00000000 ;
			12'h0000020E : data <= 8'b00000000 ;
			12'h0000020F : data <= 8'b00000000 ;
			12'h00000210 : data <= 8'b00000000 ;
			12'h00000211 : data <= 8'b00000000 ;
			12'h00000212 : data <= 8'b00011000 ;
			12'h00000213 : data <= 8'b00111100 ;
			12'h00000214 : data <= 8'b00111100 ;
			12'h00000215 : data <= 8'b00111100 ;
			12'h00000216 : data <= 8'b00011000 ;
			12'h00000217 : data <= 8'b00011000 ;
			12'h00000218 : data <= 8'b00011000 ;
			12'h00000219 : data <= 8'b00000000 ;
			12'h0000021A : data <= 8'b00011000 ;
			12'h0000021B : data <= 8'b00011000 ;
			12'h0000021C : data <= 8'b00000000 ;
			12'h0000021D : data <= 8'b00000000 ;
			12'h0000021E : data <= 8'b00000000 ;
			12'h0000021F : data <= 8'b00000000 ;
			12'h00000220 : data <= 8'b00000000 ;
			12'h00000221 : data <= 8'b01100110 ;
			12'h00000222 : data <= 8'b01100110 ;
			12'h00000223 : data <= 8'b01100110 ;
			12'h00000224 : data <= 8'b00100100 ;
			12'h00000225 : data <= 8'b00000000 ;
			12'h00000226 : data <= 8'b00000000 ;
			12'h00000227 : data <= 8'b00000000 ;
			12'h00000228 : data <= 8'b00000000 ;
			12'h00000229 : data <= 8'b00000000 ;
			12'h0000022A : data <= 8'b00000000 ;
			12'h0000022B : data <= 8'b00000000 ;
			12'h0000022C : data <= 8'b00000000 ;
			12'h0000022D : data <= 8'b00000000 ;
			12'h0000022E : data <= 8'b00000000 ;
			12'h0000022F : data <= 8'b00000000 ;
			12'h00000230 : data <= 8'b00000000 ;
			12'h00000231 : data <= 8'b00000000 ;
			12'h00000232 : data <= 8'b00000000 ;
			12'h00000233 : data <= 8'b01101100 ;
			12'h00000234 : data <= 8'b01101100 ;
			12'h00000235 : data <= 8'b11111110 ;
			12'h00000236 : data <= 8'b01101100 ;
			12'h00000237 : data <= 8'b01101100 ;
			12'h00000238 : data <= 8'b01101100 ;
			12'h00000239 : data <= 8'b11111110 ;
			12'h0000023A : data <= 8'b01101100 ;
			12'h0000023B : data <= 8'b01101100 ;
			12'h0000023C : data <= 8'b00000000 ;
			12'h0000023D : data <= 8'b00000000 ;
			12'h0000023E : data <= 8'b00000000 ;
			12'h0000023F : data <= 8'b00000000 ;
			12'h00000240 : data <= 8'b00011000 ;
			12'h00000241 : data <= 8'b00011000 ;
			12'h00000242 : data <= 8'b01111100 ;
			12'h00000243 : data <= 8'b11000110 ;
			12'h00000244 : data <= 8'b11000010 ;
			12'h00000245 : data <= 8'b11000000 ;
			12'h00000246 : data <= 8'b01111100 ;
			12'h00000247 : data <= 8'b00000110 ;
			12'h00000248 : data <= 8'b00000110 ;
			12'h00000249 : data <= 8'b10000110 ;
			12'h0000024A : data <= 8'b11000110 ;
			12'h0000024B : data <= 8'b01111100 ;
			12'h0000024C : data <= 8'b00011000 ;
			12'h0000024D : data <= 8'b00011000 ;
			12'h0000024E : data <= 8'b00000000 ;
			12'h0000024F : data <= 8'b00000000 ;
			12'h00000250 : data <= 8'b00000000 ;
			12'h00000251 : data <= 8'b00000000 ;
			12'h00000252 : data <= 8'b00000000 ;
			12'h00000253 : data <= 8'b00000000 ;
			12'h00000254 : data <= 8'b11000010 ;
			12'h00000255 : data <= 8'b11000110 ;
			12'h00000256 : data <= 8'b00001100 ;
			12'h00000257 : data <= 8'b00011000 ;
			12'h00000258 : data <= 8'b00110000 ;
			12'h00000259 : data <= 8'b01100000 ;
			12'h0000025A : data <= 8'b11000110 ;
			12'h0000025B : data <= 8'b10000110 ;
			12'h0000025C : data <= 8'b00000000 ;
			12'h0000025D : data <= 8'b00000000 ;
			12'h0000025E : data <= 8'b00000000 ;
			12'h0000025F : data <= 8'b00000000 ;
			12'h00000260 : data <= 8'b00000000 ;
			12'h00000261 : data <= 8'b00000000 ;
			12'h00000262 : data <= 8'b00111000 ;
			12'h00000263 : data <= 8'b01101100 ;
			12'h00000264 : data <= 8'b01101100 ;
			12'h00000265 : data <= 8'b00111000 ;
			12'h00000266 : data <= 8'b01110110 ;
			12'h00000267 : data <= 8'b11011100 ;
			12'h00000268 : data <= 8'b11001100 ;
			12'h00000269 : data <= 8'b11001100 ;
			12'h0000026A : data <= 8'b11001100 ;
			12'h0000026B : data <= 8'b01110110 ;
			12'h0000026C : data <= 8'b00000000 ;
			12'h0000026D : data <= 8'b00000000 ;
			12'h0000026E : data <= 8'b00000000 ;
			12'h0000026F : data <= 8'b00000000 ;
			12'h00000270 : data <= 8'b00000000 ;
			12'h00000271 : data <= 8'b00110000 ;
			12'h00000272 : data <= 8'b00110000 ;
			12'h00000273 : data <= 8'b00110000 ;
			12'h00000274 : data <= 8'b01100000 ;
			12'h00000275 : data <= 8'b00000000 ;
			12'h00000276 : data <= 8'b00000000 ;
			12'h00000277 : data <= 8'b00000000 ;
			12'h00000278 : data <= 8'b00000000 ;
			12'h00000279 : data <= 8'b00000000 ;
			12'h0000027A : data <= 8'b00000000 ;
			12'h0000027B : data <= 8'b00000000 ;
			12'h0000027C : data <= 8'b00000000 ;
			12'h0000027D : data <= 8'b00000000 ;
			12'h0000027E : data <= 8'b00000000 ;
			12'h0000027F : data <= 8'b00000000 ;
			12'h00000280 : data <= 8'b00000000 ;
			12'h00000281 : data <= 8'b00000000 ;
			12'h00000282 : data <= 8'b00001100 ;
			12'h00000283 : data <= 8'b00011000 ;
			12'h00000284 : data <= 8'b00110000 ;
			12'h00000285 : data <= 8'b00110000 ;
			12'h00000286 : data <= 8'b00110000 ;
			12'h00000287 : data <= 8'b00110000 ;
			12'h00000288 : data <= 8'b00110000 ;
			12'h00000289 : data <= 8'b00110000 ;
			12'h0000028A : data <= 8'b00011000 ;
			12'h0000028B : data <= 8'b00001100 ;
			12'h0000028C : data <= 8'b00000000 ;
			12'h0000028D : data <= 8'b00000000 ;
			12'h0000028E : data <= 8'b00000000 ;
			12'h0000028F : data <= 8'b00000000 ;
			12'h00000290 : data <= 8'b00000000 ;
			12'h00000291 : data <= 8'b00000000 ;
			12'h00000292 : data <= 8'b00110000 ;
			12'h00000293 : data <= 8'b00011000 ;
			12'h00000294 : data <= 8'b00001100 ;
			12'h00000295 : data <= 8'b00001100 ;
			12'h00000296 : data <= 8'b00001100 ;
			12'h00000297 : data <= 8'b00001100 ;
			12'h00000298 : data <= 8'b00001100 ;
			12'h00000299 : data <= 8'b00001100 ;
			12'h0000029A : data <= 8'b00011000 ;
			12'h0000029B : data <= 8'b00110000 ;
			12'h0000029C : data <= 8'b00000000 ;
			12'h0000029D : data <= 8'b00000000 ;
			12'h0000029E : data <= 8'b00000000 ;
			12'h0000029F : data <= 8'b00000000 ;
			12'h000002A0 : data <= 8'b00000000 ;
			12'h000002A1 : data <= 8'b00000000 ;
			12'h000002A2 : data <= 8'b00000000 ;
			12'h000002A3 : data <= 8'b00000000 ;
			12'h000002A4 : data <= 8'b00000000 ;
			12'h000002A5 : data <= 8'b01100110 ;
			12'h000002A6 : data <= 8'b00111100 ;
			12'h000002A7 : data <= 8'b11111111 ;
			12'h000002A8 : data <= 8'b00111100 ;
			12'h000002A9 : data <= 8'b01100110 ;
			12'h000002AA : data <= 8'b00000000 ;
			12'h000002AB : data <= 8'b00000000 ;
			12'h000002AC : data <= 8'b00000000 ;
			12'h000002AD : data <= 8'b00000000 ;
			12'h000002AE : data <= 8'b00000000 ;
			12'h000002AF : data <= 8'b00000000 ;
			12'h000002B0 : data <= 8'b00000000 ;
			12'h000002B1 : data <= 8'b00000000 ;
			12'h000002B2 : data <= 8'b00000000 ;
			12'h000002B3 : data <= 8'b00000000 ;
			12'h000002B4 : data <= 8'b00000000 ;
			12'h000002B5 : data <= 8'b00011000 ;
			12'h000002B6 : data <= 8'b00011000 ;
			12'h000002B7 : data <= 8'b01111110 ;
			12'h000002B8 : data <= 8'b00011000 ;
			12'h000002B9 : data <= 8'b00011000 ;
			12'h000002BA : data <= 8'b00000000 ;
			12'h000002BB : data <= 8'b00000000 ;
			12'h000002BC : data <= 8'b00000000 ;
			12'h000002BD : data <= 8'b00000000 ;
			12'h000002BE : data <= 8'b00000000 ;
			12'h000002BF : data <= 8'b00000000 ;
			12'h000002C0 : data <= 8'b00000000 ;
			12'h000002C1 : data <= 8'b00000000 ;
			12'h000002C2 : data <= 8'b00000000 ;
			12'h000002C3 : data <= 8'b00000000 ;
			12'h000002C4 : data <= 8'b00000000 ;
			12'h000002C5 : data <= 8'b00000000 ;
			12'h000002C6 : data <= 8'b00000000 ;
			12'h000002C7 : data <= 8'b00000000 ;
			12'h000002C8 : data <= 8'b00000000 ;
			12'h000002C9 : data <= 8'b00011000 ;
			12'h000002CA : data <= 8'b00011000 ;
			12'h000002CB : data <= 8'b00011000 ;
			12'h000002CC : data <= 8'b00110000 ;
			12'h000002CD : data <= 8'b00000000 ;
			12'h000002CE : data <= 8'b00000000 ;
			12'h000002CF : data <= 8'b00000000 ;
			12'h000002D0 : data <= 8'b00000000 ;
			12'h000002D1 : data <= 8'b00000000 ;
			12'h000002D2 : data <= 8'b00000000 ;
			12'h000002D3 : data <= 8'b00000000 ;
			12'h000002D4 : data <= 8'b00000000 ;
			12'h000002D5 : data <= 8'b00000000 ;
			12'h000002D6 : data <= 8'b00000000 ;
			12'h000002D7 : data <= 8'b11111110 ;
			12'h000002D8 : data <= 8'b00000000 ;
			12'h000002D9 : data <= 8'b00000000 ;
			12'h000002DA : data <= 8'b00000000 ;
			12'h000002DB : data <= 8'b00000000 ;
			12'h000002DC : data <= 8'b00000000 ;
			12'h000002DD : data <= 8'b00000000 ;
			12'h000002DE : data <= 8'b00000000 ;
			12'h000002DF : data <= 8'b00000000 ;
			12'h000002E0 : data <= 8'b00000000 ;
			12'h000002E1 : data <= 8'b00000000 ;
			12'h000002E2 : data <= 8'b00000000 ;
			12'h000002E3 : data <= 8'b00000000 ;
			12'h000002E4 : data <= 8'b00000000 ;
			12'h000002E5 : data <= 8'b00000000 ;
			12'h000002E6 : data <= 8'b00000000 ;
			12'h000002E7 : data <= 8'b00000000 ;
			12'h000002E8 : data <= 8'b00000000 ;
			12'h000002E9 : data <= 8'b00000000 ;
			12'h000002EA : data <= 8'b00011000 ;
			12'h000002EB : data <= 8'b00011000 ;
			12'h000002EC : data <= 8'b00000000 ;
			12'h000002ED : data <= 8'b00000000 ;
			12'h000002EE : data <= 8'b00000000 ;
			12'h000002EF : data <= 8'b00000000 ;
			12'h000002F0 : data <= 8'b00000000 ;
			12'h000002F1 : data <= 8'b00000000 ;
			12'h000002F2 : data <= 8'b00000000 ;
			12'h000002F3 : data <= 8'b00000000 ;
			12'h000002F4 : data <= 8'b00000010 ;
			12'h000002F5 : data <= 8'b00000110 ;
			12'h000002F6 : data <= 8'b00001100 ;
			12'h000002F7 : data <= 8'b00011000 ;
			12'h000002F8 : data <= 8'b00110000 ;
			12'h000002F9 : data <= 8'b01100000 ;
			12'h000002FA : data <= 8'b11000000 ;
			12'h000002FB : data <= 8'b10000000 ;
			12'h000002FC : data <= 8'b00000000 ;
			12'h000002FD : data <= 8'b00000000 ;
			12'h000002FE : data <= 8'b00000000 ;
			12'h000002FF : data <= 8'b00000000 ;
			12'h00000300 : data <= 8'b00000000 ;
			12'h00000301 : data <= 8'b00000000 ;
			12'h00000302 : data <= 8'b00111000 ;
			12'h00000303 : data <= 8'b01101100 ;
			12'h00000304 : data <= 8'b11000110 ;
			12'h00000305 : data <= 8'b11000110 ;
			12'h00000306 : data <= 8'b11010110 ;
			12'h00000307 : data <= 8'b11010110 ;
			12'h00000308 : data <= 8'b11000110 ;
			12'h00000309 : data <= 8'b11000110 ;
			12'h0000030A : data <= 8'b01101100 ;
			12'h0000030B : data <= 8'b00111000 ;
			12'h0000030C : data <= 8'b00000000 ;
			12'h0000030D : data <= 8'b00000000 ;
			12'h0000030E : data <= 8'b00000000 ;
			12'h0000030F : data <= 8'b00000000 ;
			12'h00000310 : data <= 8'b00000000 ;
			12'h00000311 : data <= 8'b00000000 ;
			12'h00000312 : data <= 8'b00011000 ;
			12'h00000313 : data <= 8'b00111000 ;
			12'h00000314 : data <= 8'b01111000 ;
			12'h00000315 : data <= 8'b00011000 ;
			12'h00000316 : data <= 8'b00011000 ;
			12'h00000317 : data <= 8'b00011000 ;
			12'h00000318 : data <= 8'b00011000 ;
			12'h00000319 : data <= 8'b00011000 ;
			12'h0000031A : data <= 8'b00011000 ;
			12'h0000031B : data <= 8'b01111110 ;
			12'h0000031C : data <= 8'b00000000 ;
			12'h0000031D : data <= 8'b00000000 ;
			12'h0000031E : data <= 8'b00000000 ;
			12'h0000031F : data <= 8'b00000000 ;
			12'h00000320 : data <= 8'b00000000 ;
			12'h00000321 : data <= 8'b00000000 ;
			12'h00000322 : data <= 8'b01111100 ;
			12'h00000323 : data <= 8'b11000110 ;
			12'h00000324 : data <= 8'b00000110 ;
			12'h00000325 : data <= 8'b00001100 ;
			12'h00000326 : data <= 8'b00011000 ;
			12'h00000327 : data <= 8'b00110000 ;
			12'h00000328 : data <= 8'b01100000 ;
			12'h00000329 : data <= 8'b11000000 ;
			12'h0000032A : data <= 8'b11000110 ;
			12'h0000032B : data <= 8'b11111110 ;
			12'h0000032C : data <= 8'b00000000 ;
			12'h0000032D : data <= 8'b00000000 ;
			12'h0000032E : data <= 8'b00000000 ;
			12'h0000032F : data <= 8'b00000000 ;
			12'h00000330 : data <= 8'b00000000 ;
			12'h00000331 : data <= 8'b00000000 ;
			12'h00000332 : data <= 8'b01111100 ;
			12'h00000333 : data <= 8'b11000110 ;
			12'h00000334 : data <= 8'b00000110 ;
			12'h00000335 : data <= 8'b00000110 ;
			12'h00000336 : data <= 8'b00111100 ;
			12'h00000337 : data <= 8'b00000110 ;
			12'h00000338 : data <= 8'b00000110 ;
			12'h00000339 : data <= 8'b00000110 ;
			12'h0000033A : data <= 8'b11000110 ;
			12'h0000033B : data <= 8'b01111100 ;
			12'h0000033C : data <= 8'b00000000 ;
			12'h0000033D : data <= 8'b00000000 ;
			12'h0000033E : data <= 8'b00000000 ;
			12'h0000033F : data <= 8'b00000000 ;
			12'h00000340 : data <= 8'b00000000 ;
			12'h00000341 : data <= 8'b00000000 ;
			12'h00000342 : data <= 8'b00001100 ;
			12'h00000343 : data <= 8'b00011100 ;
			12'h00000344 : data <= 8'b00111100 ;
			12'h00000345 : data <= 8'b01101100 ;
			12'h00000346 : data <= 8'b11001100 ;
			12'h00000347 : data <= 8'b11111110 ;
			12'h00000348 : data <= 8'b00001100 ;
			12'h00000349 : data <= 8'b00001100 ;
			12'h0000034A : data <= 8'b00001100 ;
			12'h0000034B : data <= 8'b00011110 ;
			12'h0000034C : data <= 8'b00000000 ;
			12'h0000034D : data <= 8'b00000000 ;
			12'h0000034E : data <= 8'b00000000 ;
			12'h0000034F : data <= 8'b00000000 ;
			12'h00000350 : data <= 8'b00000000 ;
			12'h00000351 : data <= 8'b00000000 ;
			12'h00000352 : data <= 8'b11111110 ;
			12'h00000353 : data <= 8'b11000000 ;
			12'h00000354 : data <= 8'b11000000 ;
			12'h00000355 : data <= 8'b11000000 ;
			12'h00000356 : data <= 8'b11111100 ;
			12'h00000357 : data <= 8'b00000110 ;
			12'h00000358 : data <= 8'b00000110 ;
			12'h00000359 : data <= 8'b00000110 ;
			12'h0000035A : data <= 8'b11000110 ;
			12'h0000035B : data <= 8'b01111100 ;
			12'h0000035C : data <= 8'b00000000 ;
			12'h0000035D : data <= 8'b00000000 ;
			12'h0000035E : data <= 8'b00000000 ;
			12'h0000035F : data <= 8'b00000000 ;
			12'h00000360 : data <= 8'b00000000 ;
			12'h00000361 : data <= 8'b00000000 ;
			12'h00000362 : data <= 8'b00111000 ;
			12'h00000363 : data <= 8'b01100000 ;
			12'h00000364 : data <= 8'b11000000 ;
			12'h00000365 : data <= 8'b11000000 ;
			12'h00000366 : data <= 8'b11111100 ;
			12'h00000367 : data <= 8'b11000110 ;
			12'h00000368 : data <= 8'b11000110 ;
			12'h00000369 : data <= 8'b11000110 ;
			12'h0000036A : data <= 8'b11000110 ;
			12'h0000036B : data <= 8'b01111100 ;
			12'h0000036C : data <= 8'b00000000 ;
			12'h0000036D : data <= 8'b00000000 ;
			12'h0000036E : data <= 8'b00000000 ;
			12'h0000036F : data <= 8'b00000000 ;
			12'h00000370 : data <= 8'b00000000 ;
			12'h00000371 : data <= 8'b00000000 ;
			12'h00000372 : data <= 8'b11111110 ;
			12'h00000373 : data <= 8'b11000110 ;
			12'h00000374 : data <= 8'b00000110 ;
			12'h00000375 : data <= 8'b00000110 ;
			12'h00000376 : data <= 8'b00001100 ;
			12'h00000377 : data <= 8'b00011000 ;
			12'h00000378 : data <= 8'b00110000 ;
			12'h00000379 : data <= 8'b00110000 ;
			12'h0000037A : data <= 8'b00110000 ;
			12'h0000037B : data <= 8'b00110000 ;
			12'h0000037C : data <= 8'b00000000 ;
			12'h0000037D : data <= 8'b00000000 ;
			12'h0000037E : data <= 8'b00000000 ;
			12'h0000037F : data <= 8'b00000000 ;
			12'h00000380 : data <= 8'b00000000 ;
			12'h00000381 : data <= 8'b00000000 ;
			12'h00000382 : data <= 8'b01111100 ;
			12'h00000383 : data <= 8'b11000110 ;
			12'h00000384 : data <= 8'b11000110 ;
			12'h00000385 : data <= 8'b11000110 ;
			12'h00000386 : data <= 8'b01111100 ;
			12'h00000387 : data <= 8'b11000110 ;
			12'h00000388 : data <= 8'b11000110 ;
			12'h00000389 : data <= 8'b11000110 ;
			12'h0000038A : data <= 8'b11000110 ;
			12'h0000038B : data <= 8'b01111100 ;
			12'h0000038C : data <= 8'b00000000 ;
			12'h0000038D : data <= 8'b00000000 ;
			12'h0000038E : data <= 8'b00000000 ;
			12'h0000038F : data <= 8'b00000000 ;
			12'h00000390 : data <= 8'b00000000 ;
			12'h00000391 : data <= 8'b00000000 ;
			12'h00000392 : data <= 8'b01111100 ;
			12'h00000393 : data <= 8'b11000110 ;
			12'h00000394 : data <= 8'b11000110 ;
			12'h00000395 : data <= 8'b11000110 ;
			12'h00000396 : data <= 8'b01111110 ;
			12'h00000397 : data <= 8'b00000110 ;
			12'h00000398 : data <= 8'b00000110 ;
			12'h00000399 : data <= 8'b00000110 ;
			12'h0000039A : data <= 8'b00001100 ;
			12'h0000039B : data <= 8'b01111000 ;
			12'h0000039C : data <= 8'b00000000 ;
			12'h0000039D : data <= 8'b00000000 ;
			12'h0000039E : data <= 8'b00000000 ;
			12'h0000039F : data <= 8'b00000000 ;
			12'h000003A0 : data <= 8'b00000000 ;
			12'h000003A1 : data <= 8'b00000000 ;
			12'h000003A2 : data <= 8'b00000000 ;
			12'h000003A3 : data <= 8'b00000000 ;
			12'h000003A4 : data <= 8'b00011000 ;
			12'h000003A5 : data <= 8'b00011000 ;
			12'h000003A6 : data <= 8'b00000000 ;
			12'h000003A7 : data <= 8'b00000000 ;
			12'h000003A8 : data <= 8'b00000000 ;
			12'h000003A9 : data <= 8'b00011000 ;
			12'h000003AA : data <= 8'b00011000 ;
			12'h000003AB : data <= 8'b00000000 ;
			12'h000003AC : data <= 8'b00000000 ;
			12'h000003AD : data <= 8'b00000000 ;
			12'h000003AE : data <= 8'b00000000 ;
			12'h000003AF : data <= 8'b00000000 ;
			12'h000003B0 : data <= 8'b00000000 ;
			12'h000003B1 : data <= 8'b00000000 ;
			12'h000003B2 : data <= 8'b00000000 ;
			12'h000003B3 : data <= 8'b00000000 ;
			12'h000003B4 : data <= 8'b00011000 ;
			12'h000003B5 : data <= 8'b00011000 ;
			12'h000003B6 : data <= 8'b00000000 ;
			12'h000003B7 : data <= 8'b00000000 ;
			12'h000003B8 : data <= 8'b00000000 ;
			12'h000003B9 : data <= 8'b00011000 ;
			12'h000003BA : data <= 8'b00011000 ;
			12'h000003BB : data <= 8'b00110000 ;
			12'h000003BC : data <= 8'b00000000 ;
			12'h000003BD : data <= 8'b00000000 ;
			12'h000003BE : data <= 8'b00000000 ;
			12'h000003BF : data <= 8'b00000000 ;
			12'h000003C0 : data <= 8'b00000000 ;
			12'h000003C1 : data <= 8'b00000000 ;
			12'h000003C2 : data <= 8'b00000000 ;
			12'h000003C3 : data <= 8'b00000110 ;
			12'h000003C4 : data <= 8'b00001100 ;
			12'h000003C5 : data <= 8'b00011000 ;
			12'h000003C6 : data <= 8'b00110000 ;
			12'h000003C7 : data <= 8'b01100000 ;
			12'h000003C8 : data <= 8'b00110000 ;
			12'h000003C9 : data <= 8'b00011000 ;
			12'h000003CA : data <= 8'b00001100 ;
			12'h000003CB : data <= 8'b00000110 ;
			12'h000003CC : data <= 8'b00000000 ;
			12'h000003CD : data <= 8'b00000000 ;
			12'h000003CE : data <= 8'b00000000 ;
			12'h000003CF : data <= 8'b00000000 ;
			12'h000003D0 : data <= 8'b00000000 ;
			12'h000003D1 : data <= 8'b00000000 ;
			12'h000003D2 : data <= 8'b00000000 ;
			12'h000003D3 : data <= 8'b00000000 ;
			12'h000003D4 : data <= 8'b00000000 ;
			12'h000003D5 : data <= 8'b01111110 ;
			12'h000003D6 : data <= 8'b00000000 ;
			12'h000003D7 : data <= 8'b00000000 ;
			12'h000003D8 : data <= 8'b01111110 ;
			12'h000003D9 : data <= 8'b00000000 ;
			12'h000003DA : data <= 8'b00000000 ;
			12'h000003DB : data <= 8'b00000000 ;
			12'h000003DC : data <= 8'b00000000 ;
			12'h000003DD : data <= 8'b00000000 ;
			12'h000003DE : data <= 8'b00000000 ;
			12'h000003DF : data <= 8'b00000000 ;
			12'h000003E0 : data <= 8'b00000000 ;
			12'h000003E1 : data <= 8'b00000000 ;
			12'h000003E2 : data <= 8'b00000000 ;
			12'h000003E3 : data <= 8'b01100000 ;
			12'h000003E4 : data <= 8'b00110000 ;
			12'h000003E5 : data <= 8'b00011000 ;
			12'h000003E6 : data <= 8'b00001100 ;
			12'h000003E7 : data <= 8'b00000110 ;
			12'h000003E8 : data <= 8'b00001100 ;
			12'h000003E9 : data <= 8'b00011000 ;
			12'h000003EA : data <= 8'b00110000 ;
			12'h000003EB : data <= 8'b01100000 ;
			12'h000003EC : data <= 8'b00000000 ;
			12'h000003ED : data <= 8'b00000000 ;
			12'h000003EE : data <= 8'b00000000 ;
			12'h000003EF : data <= 8'b00000000 ;
			12'h000003F0 : data <= 8'b00000000 ;
			12'h000003F1 : data <= 8'b00000000 ;
			12'h000003F2 : data <= 8'b01111100 ;
			12'h000003F3 : data <= 8'b11000110 ;
			12'h000003F4 : data <= 8'b11000110 ;
			12'h000003F5 : data <= 8'b00001100 ;
			12'h000003F6 : data <= 8'b00011000 ;
			12'h000003F7 : data <= 8'b00011000 ;
			12'h000003F8 : data <= 8'b00011000 ;
			12'h000003F9 : data <= 8'b00000000 ;
			12'h000003FA : data <= 8'b00011000 ;
			12'h000003FB : data <= 8'b00011000 ;
			12'h000003FC : data <= 8'b00000000 ;
			12'h000003FD : data <= 8'b00000000 ;
			12'h000003FE : data <= 8'b00000000 ;
			12'h000003FF : data <= 8'b00000000 ;
			12'h00000400 : data <= 8'b00000000 ;
			12'h00000401 : data <= 8'b00000000 ;
			12'h00000402 : data <= 8'b00000000 ;
			12'h00000403 : data <= 8'b01111100 ;
			12'h00000404 : data <= 8'b11000110 ;
			12'h00000405 : data <= 8'b11000110 ;
			12'h00000406 : data <= 8'b11011110 ;
			12'h00000407 : data <= 8'b11011110 ;
			12'h00000408 : data <= 8'b11011110 ;
			12'h00000409 : data <= 8'b11011100 ;
			12'h0000040A : data <= 8'b11000000 ;
			12'h0000040B : data <= 8'b01111100 ;
			12'h0000040C : data <= 8'b00000000 ;
			12'h0000040D : data <= 8'b00000000 ;
			12'h0000040E : data <= 8'b00000000 ;
			12'h0000040F : data <= 8'b00000000 ;
			12'h00000410 : data <= 8'b00000000 ;
			12'h00000411 : data <= 8'b00000000 ;
			12'h00000412 : data <= 8'b00010000 ;
			12'h00000413 : data <= 8'b00111000 ;
			12'h00000414 : data <= 8'b01101100 ;
			12'h00000415 : data <= 8'b11000110 ;
			12'h00000416 : data <= 8'b11000110 ;
			12'h00000417 : data <= 8'b11111110 ;
			12'h00000418 : data <= 8'b11000110 ;
			12'h00000419 : data <= 8'b11000110 ;
			12'h0000041A : data <= 8'b11000110 ;
			12'h0000041B : data <= 8'b11000110 ;
			12'h0000041C : data <= 8'b00000000 ;
			12'h0000041D : data <= 8'b00000000 ;
			12'h0000041E : data <= 8'b00000000 ;
			12'h0000041F : data <= 8'b00000000 ;
			12'h00000420 : data <= 8'b00000000 ;
			12'h00000421 : data <= 8'b00000000 ;
			12'h00000422 : data <= 8'b11111100 ;
			12'h00000423 : data <= 8'b01100110 ;
			12'h00000424 : data <= 8'b01100110 ;
			12'h00000425 : data <= 8'b01100110 ;
			12'h00000426 : data <= 8'b01111100 ;
			12'h00000427 : data <= 8'b01100110 ;
			12'h00000428 : data <= 8'b01100110 ;
			12'h00000429 : data <= 8'b01100110 ;
			12'h0000042A : data <= 8'b01100110 ;
			12'h0000042B : data <= 8'b11111100 ;
			12'h0000042C : data <= 8'b00000000 ;
			12'h0000042D : data <= 8'b00000000 ;
			12'h0000042E : data <= 8'b00000000 ;
			12'h0000042F : data <= 8'b00000000 ;
			12'h00000430 : data <= 8'b00000000 ;
			12'h00000431 : data <= 8'b00000000 ;
			12'h00000432 : data <= 8'b00111100 ;
			12'h00000433 : data <= 8'b01100110 ;
			12'h00000434 : data <= 8'b11000010 ;
			12'h00000435 : data <= 8'b11000000 ;
			12'h00000436 : data <= 8'b11000000 ;
			12'h00000437 : data <= 8'b11000000 ;
			12'h00000438 : data <= 8'b11000000 ;
			12'h00000439 : data <= 8'b11000010 ;
			12'h0000043A : data <= 8'b01100110 ;
			12'h0000043B : data <= 8'b00111100 ;
			12'h0000043C : data <= 8'b00000000 ;
			12'h0000043D : data <= 8'b00000000 ;
			12'h0000043E : data <= 8'b00000000 ;
			12'h0000043F : data <= 8'b00000000 ;
			12'h00000440 : data <= 8'b00000000 ;
			12'h00000441 : data <= 8'b00000000 ;
			12'h00000442 : data <= 8'b11111000 ;
			12'h00000443 : data <= 8'b01101100 ;
			12'h00000444 : data <= 8'b01100110 ;
			12'h00000445 : data <= 8'b01100110 ;
			12'h00000446 : data <= 8'b01100110 ;
			12'h00000447 : data <= 8'b01100110 ;
			12'h00000448 : data <= 8'b01100110 ;
			12'h00000449 : data <= 8'b01100110 ;
			12'h0000044A : data <= 8'b01101100 ;
			12'h0000044B : data <= 8'b11111000 ;
			12'h0000044C : data <= 8'b00000000 ;
			12'h0000044D : data <= 8'b00000000 ;
			12'h0000044E : data <= 8'b00000000 ;
			12'h0000044F : data <= 8'b00000000 ;
			12'h00000450 : data <= 8'b00000000 ;
			12'h00000451 : data <= 8'b00000000 ;
			12'h00000452 : data <= 8'b11111110 ;
			12'h00000453 : data <= 8'b01100110 ;
			12'h00000454 : data <= 8'b01100010 ;
			12'h00000455 : data <= 8'b01101000 ;
			12'h00000456 : data <= 8'b01111000 ;
			12'h00000457 : data <= 8'b01101000 ;
			12'h00000458 : data <= 8'b01100000 ;
			12'h00000459 : data <= 8'b01100010 ;
			12'h0000045A : data <= 8'b01100110 ;
			12'h0000045B : data <= 8'b11111110 ;
			12'h0000045C : data <= 8'b00000000 ;
			12'h0000045D : data <= 8'b00000000 ;
			12'h0000045E : data <= 8'b00000000 ;
			12'h0000045F : data <= 8'b00000000 ;
			12'h00000460 : data <= 8'b00000000 ;
			12'h00000461 : data <= 8'b00000000 ;
			12'h00000462 : data <= 8'b11111110 ;
			12'h00000463 : data <= 8'b01100110 ;
			12'h00000464 : data <= 8'b01100010 ;
			12'h00000465 : data <= 8'b01101000 ;
			12'h00000466 : data <= 8'b01111000 ;
			12'h00000467 : data <= 8'b01101000 ;
			12'h00000468 : data <= 8'b01100000 ;
			12'h00000469 : data <= 8'b01100000 ;
			12'h0000046A : data <= 8'b01100000 ;
			12'h0000046B : data <= 8'b11110000 ;
			12'h0000046C : data <= 8'b00000000 ;
			12'h0000046D : data <= 8'b00000000 ;
			12'h0000046E : data <= 8'b00000000 ;
			12'h0000046F : data <= 8'b00000000 ;
			12'h00000470 : data <= 8'b00000000 ;
			12'h00000471 : data <= 8'b00000000 ;
			12'h00000472 : data <= 8'b00111100 ;
			12'h00000473 : data <= 8'b01100110 ;
			12'h00000474 : data <= 8'b11000010 ;
			12'h00000475 : data <= 8'b11000000 ;
			12'h00000476 : data <= 8'b11000000 ;
			12'h00000477 : data <= 8'b11011110 ;
			12'h00000478 : data <= 8'b11000110 ;
			12'h00000479 : data <= 8'b11000110 ;
			12'h0000047A : data <= 8'b01100110 ;
			12'h0000047B : data <= 8'b00111010 ;
			12'h0000047C : data <= 8'b00000000 ;
			12'h0000047D : data <= 8'b00000000 ;
			12'h0000047E : data <= 8'b00000000 ;
			12'h0000047F : data <= 8'b00000000 ;
			12'h00000480 : data <= 8'b00000000 ;
			12'h00000481 : data <= 8'b00000000 ;
			12'h00000482 : data <= 8'b11000110 ;
			12'h00000483 : data <= 8'b11000110 ;
			12'h00000484 : data <= 8'b11000110 ;
			12'h00000485 : data <= 8'b11000110 ;
			12'h00000486 : data <= 8'b11111110 ;
			12'h00000487 : data <= 8'b11000110 ;
			12'h00000488 : data <= 8'b11000110 ;
			12'h00000489 : data <= 8'b11000110 ;
			12'h0000048A : data <= 8'b11000110 ;
			12'h0000048B : data <= 8'b11000110 ;
			12'h0000048C : data <= 8'b00000000 ;
			12'h0000048D : data <= 8'b00000000 ;
			12'h0000048E : data <= 8'b00000000 ;
			12'h0000048F : data <= 8'b00000000 ;
			12'h00000490 : data <= 8'b00000000 ;
			12'h00000491 : data <= 8'b00000000 ;
			12'h00000492 : data <= 8'b00111100 ;
			12'h00000493 : data <= 8'b00011000 ;
			12'h00000494 : data <= 8'b00011000 ;
			12'h00000495 : data <= 8'b00011000 ;
			12'h00000496 : data <= 8'b00011000 ;
			12'h00000497 : data <= 8'b00011000 ;
			12'h00000498 : data <= 8'b00011000 ;
			12'h00000499 : data <= 8'b00011000 ;
			12'h0000049A : data <= 8'b00011000 ;
			12'h0000049B : data <= 8'b00111100 ;
			12'h0000049C : data <= 8'b00000000 ;
			12'h0000049D : data <= 8'b00000000 ;
			12'h0000049E : data <= 8'b00000000 ;
			12'h0000049F : data <= 8'b00000000 ;
			12'h000004A0 : data <= 8'b00000000 ;
			12'h000004A1 : data <= 8'b00000000 ;
			12'h000004A2 : data <= 8'b00011110 ;
			12'h000004A3 : data <= 8'b00001100 ;
			12'h000004A4 : data <= 8'b00001100 ;
			12'h000004A5 : data <= 8'b00001100 ;
			12'h000004A6 : data <= 8'b00001100 ;
			12'h000004A7 : data <= 8'b00001100 ;
			12'h000004A8 : data <= 8'b11001100 ;
			12'h000004A9 : data <= 8'b11001100 ;
			12'h000004AA : data <= 8'b11001100 ;
			12'h000004AB : data <= 8'b01111000 ;
			12'h000004AC : data <= 8'b00000000 ;
			12'h000004AD : data <= 8'b00000000 ;
			12'h000004AE : data <= 8'b00000000 ;
			12'h000004AF : data <= 8'b00000000 ;
			12'h000004B0 : data <= 8'b00000000 ;
			12'h000004B1 : data <= 8'b00000000 ;
			12'h000004B2 : data <= 8'b11100110 ;
			12'h000004B3 : data <= 8'b01100110 ;
			12'h000004B4 : data <= 8'b01100110 ;
			12'h000004B5 : data <= 8'b01101100 ;
			12'h000004B6 : data <= 8'b01111000 ;
			12'h000004B7 : data <= 8'b01111000 ;
			12'h000004B8 : data <= 8'b01101100 ;
			12'h000004B9 : data <= 8'b01100110 ;
			12'h000004BA : data <= 8'b01100110 ;
			12'h000004BB : data <= 8'b11100110 ;
			12'h000004BC : data <= 8'b00000000 ;
			12'h000004BD : data <= 8'b00000000 ;
			12'h000004BE : data <= 8'b00000000 ;
			12'h000004BF : data <= 8'b00000000 ;
			12'h000004C0 : data <= 8'b00000000 ;
			12'h000004C1 : data <= 8'b00000000 ;
			12'h000004C2 : data <= 8'b11110000 ;
			12'h000004C3 : data <= 8'b01100000 ;
			12'h000004C4 : data <= 8'b01100000 ;
			12'h000004C5 : data <= 8'b01100000 ;
			12'h000004C6 : data <= 8'b01100000 ;
			12'h000004C7 : data <= 8'b01100000 ;
			12'h000004C8 : data <= 8'b01100000 ;
			12'h000004C9 : data <= 8'b01100010 ;
			12'h000004CA : data <= 8'b01100110 ;
			12'h000004CB : data <= 8'b11111110 ;
			12'h000004CC : data <= 8'b00000000 ;
			12'h000004CD : data <= 8'b00000000 ;
			12'h000004CE : data <= 8'b00000000 ;
			12'h000004CF : data <= 8'b00000000 ;
			12'h000004D0 : data <= 8'b00000000 ;
			12'h000004D1 : data <= 8'b00000000 ;
			12'h000004D2 : data <= 8'b11000110 ;
			12'h000004D3 : data <= 8'b11101110 ;
			12'h000004D4 : data <= 8'b11111110 ;
			12'h000004D5 : data <= 8'b11111110 ;
			12'h000004D6 : data <= 8'b11010110 ;
			12'h000004D7 : data <= 8'b11000110 ;
			12'h000004D8 : data <= 8'b11000110 ;
			12'h000004D9 : data <= 8'b11000110 ;
			12'h000004DA : data <= 8'b11000110 ;
			12'h000004DB : data <= 8'b11000110 ;
			12'h000004DC : data <= 8'b00000000 ;
			12'h000004DD : data <= 8'b00000000 ;
			12'h000004DE : data <= 8'b00000000 ;
			12'h000004DF : data <= 8'b00000000 ;
			12'h000004E0 : data <= 8'b00000000 ;
			12'h000004E1 : data <= 8'b00000000 ;
			12'h000004E2 : data <= 8'b11000110 ;
			12'h000004E3 : data <= 8'b11100110 ;
			12'h000004E4 : data <= 8'b11110110 ;
			12'h000004E5 : data <= 8'b11111110 ;
			12'h000004E6 : data <= 8'b11011110 ;
			12'h000004E7 : data <= 8'b11001110 ;
			12'h000004E8 : data <= 8'b11000110 ;
			12'h000004E9 : data <= 8'b11000110 ;
			12'h000004EA : data <= 8'b11000110 ;
			12'h000004EB : data <= 8'b11000110 ;
			12'h000004EC : data <= 8'b00000000 ;
			12'h000004ED : data <= 8'b00000000 ;
			12'h000004EE : data <= 8'b00000000 ;
			12'h000004EF : data <= 8'b00000000 ;
			12'h000004F0 : data <= 8'b00000000 ;
			12'h000004F1 : data <= 8'b00000000 ;
			12'h000004F2 : data <= 8'b01111100 ;
			12'h000004F3 : data <= 8'b11000110 ;
			12'h000004F4 : data <= 8'b11000110 ;
			12'h000004F5 : data <= 8'b11000110 ;
			12'h000004F6 : data <= 8'b11000110 ;
			12'h000004F7 : data <= 8'b11000110 ;
			12'h000004F8 : data <= 8'b11000110 ;
			12'h000004F9 : data <= 8'b11000110 ;
			12'h000004FA : data <= 8'b11000110 ;
			12'h000004FB : data <= 8'b01111100 ;
			12'h000004FC : data <= 8'b00000000 ;
			12'h000004FD : data <= 8'b00000000 ;
			12'h000004FE : data <= 8'b00000000 ;
			12'h000004FF : data <= 8'b00000000 ;
			12'h00000500 : data <= 8'b00000000 ;
			12'h00000501 : data <= 8'b00000000 ;
			12'h00000502 : data <= 8'b11111100 ;
			12'h00000503 : data <= 8'b01100110 ;
			12'h00000504 : data <= 8'b01100110 ;
			12'h00000505 : data <= 8'b01100110 ;
			12'h00000506 : data <= 8'b01111100 ;
			12'h00000507 : data <= 8'b01100000 ;
			12'h00000508 : data <= 8'b01100000 ;
			12'h00000509 : data <= 8'b01100000 ;
			12'h0000050A : data <= 8'b01100000 ;
			12'h0000050B : data <= 8'b11110000 ;
			12'h0000050C : data <= 8'b00000000 ;
			12'h0000050D : data <= 8'b00000000 ;
			12'h0000050E : data <= 8'b00000000 ;
			12'h0000050F : data <= 8'b00000000 ;
			12'h00000510 : data <= 8'b00000000 ;
			12'h00000511 : data <= 8'b00000000 ;
			12'h00000512 : data <= 8'b01111100 ;
			12'h00000513 : data <= 8'b11000110 ;
			12'h00000514 : data <= 8'b11000110 ;
			12'h00000515 : data <= 8'b11000110 ;
			12'h00000516 : data <= 8'b11000110 ;
			12'h00000517 : data <= 8'b11000110 ;
			12'h00000518 : data <= 8'b11000110 ;
			12'h00000519 : data <= 8'b11010110 ;
			12'h0000051A : data <= 8'b11011110 ;
			12'h0000051B : data <= 8'b01111100 ;
			12'h0000051C : data <= 8'b00001100 ;
			12'h0000051D : data <= 8'b00001110 ;
			12'h0000051E : data <= 8'b00000000 ;
			12'h0000051F : data <= 8'b00000000 ;
			12'h00000520 : data <= 8'b00000000 ;
			12'h00000521 : data <= 8'b00000000 ;
			12'h00000522 : data <= 8'b11111100 ;
			12'h00000523 : data <= 8'b01100110 ;
			12'h00000524 : data <= 8'b01100110 ;
			12'h00000525 : data <= 8'b01100110 ;
			12'h00000526 : data <= 8'b01111100 ;
			12'h00000527 : data <= 8'b01101100 ;
			12'h00000528 : data <= 8'b01100110 ;
			12'h00000529 : data <= 8'b01100110 ;
			12'h0000052A : data <= 8'b01100110 ;
			12'h0000052B : data <= 8'b11100110 ;
			12'h0000052C : data <= 8'b00000000 ;
			12'h0000052D : data <= 8'b00000000 ;
			12'h0000052E : data <= 8'b00000000 ;
			12'h0000052F : data <= 8'b00000000 ;
			12'h00000530 : data <= 8'b00000000 ;
			12'h00000531 : data <= 8'b00000000 ;
			12'h00000532 : data <= 8'b01111100 ;
			12'h00000533 : data <= 8'b11000110 ;
			12'h00000534 : data <= 8'b11000110 ;
			12'h00000535 : data <= 8'b01100000 ;
			12'h00000536 : data <= 8'b00111000 ;
			12'h00000537 : data <= 8'b00001100 ;
			12'h00000538 : data <= 8'b00000110 ;
			12'h00000539 : data <= 8'b11000110 ;
			12'h0000053A : data <= 8'b11000110 ;
			12'h0000053B : data <= 8'b01111100 ;
			12'h0000053C : data <= 8'b00000000 ;
			12'h0000053D : data <= 8'b00000000 ;
			12'h0000053E : data <= 8'b00000000 ;
			12'h0000053F : data <= 8'b00000000 ;
			12'h00000540 : data <= 8'b00000000 ;
			12'h00000541 : data <= 8'b00000000 ;
			12'h00000542 : data <= 8'b01111110 ;
			12'h00000543 : data <= 8'b01111110 ;
			12'h00000544 : data <= 8'b01011010 ;
			12'h00000545 : data <= 8'b00011000 ;
			12'h00000546 : data <= 8'b00011000 ;
			12'h00000547 : data <= 8'b00011000 ;
			12'h00000548 : data <= 8'b00011000 ;
			12'h00000549 : data <= 8'b00011000 ;
			12'h0000054A : data <= 8'b00011000 ;
			12'h0000054B : data <= 8'b00111100 ;
			12'h0000054C : data <= 8'b00000000 ;
			12'h0000054D : data <= 8'b00000000 ;
			12'h0000054E : data <= 8'b00000000 ;
			12'h0000054F : data <= 8'b00000000 ;
			12'h00000550 : data <= 8'b00000000 ;
			12'h00000551 : data <= 8'b00000000 ;
			12'h00000552 : data <= 8'b11000110 ;
			12'h00000553 : data <= 8'b11000110 ;
			12'h00000554 : data <= 8'b11000110 ;
			12'h00000555 : data <= 8'b11000110 ;
			12'h00000556 : data <= 8'b11000110 ;
			12'h00000557 : data <= 8'b11000110 ;
			12'h00000558 : data <= 8'b11000110 ;
			12'h00000559 : data <= 8'b11000110 ;
			12'h0000055A : data <= 8'b11000110 ;
			12'h0000055B : data <= 8'b01111100 ;
			12'h0000055C : data <= 8'b00000000 ;
			12'h0000055D : data <= 8'b00000000 ;
			12'h0000055E : data <= 8'b00000000 ;
			12'h0000055F : data <= 8'b00000000 ;
			12'h00000560 : data <= 8'b00000000 ;
			12'h00000561 : data <= 8'b00000000 ;
			12'h00000562 : data <= 8'b11000110 ;
			12'h00000563 : data <= 8'b11000110 ;
			12'h00000564 : data <= 8'b11000110 ;
			12'h00000565 : data <= 8'b11000110 ;
			12'h00000566 : data <= 8'b11000110 ;
			12'h00000567 : data <= 8'b11000110 ;
			12'h00000568 : data <= 8'b11000110 ;
			12'h00000569 : data <= 8'b01101100 ;
			12'h0000056A : data <= 8'b00111000 ;
			12'h0000056B : data <= 8'b00010000 ;
			12'h0000056C : data <= 8'b00000000 ;
			12'h0000056D : data <= 8'b00000000 ;
			12'h0000056E : data <= 8'b00000000 ;
			12'h0000056F : data <= 8'b00000000 ;
			12'h00000570 : data <= 8'b00000000 ;
			12'h00000571 : data <= 8'b00000000 ;
			12'h00000572 : data <= 8'b11000110 ;
			12'h00000573 : data <= 8'b11000110 ;
			12'h00000574 : data <= 8'b11000110 ;
			12'h00000575 : data <= 8'b11000110 ;
			12'h00000576 : data <= 8'b11010110 ;
			12'h00000577 : data <= 8'b11010110 ;
			12'h00000578 : data <= 8'b11010110 ;
			12'h00000579 : data <= 8'b11111110 ;
			12'h0000057A : data <= 8'b11101110 ;
			12'h0000057B : data <= 8'b01101100 ;
			12'h0000057C : data <= 8'b00000000 ;
			12'h0000057D : data <= 8'b00000000 ;
			12'h0000057E : data <= 8'b00000000 ;
			12'h0000057F : data <= 8'b00000000 ;
			12'h00000580 : data <= 8'b00000000 ;
			12'h00000581 : data <= 8'b00000000 ;
			12'h00000582 : data <= 8'b11000110 ;
			12'h00000583 : data <= 8'b11000110 ;
			12'h00000584 : data <= 8'b01101100 ;
			12'h00000585 : data <= 8'b01111100 ;
			12'h00000586 : data <= 8'b00111000 ;
			12'h00000587 : data <= 8'b00111000 ;
			12'h00000588 : data <= 8'b01111100 ;
			12'h00000589 : data <= 8'b01101100 ;
			12'h0000058A : data <= 8'b11000110 ;
			12'h0000058B : data <= 8'b11000110 ;
			12'h0000058C : data <= 8'b00000000 ;
			12'h0000058D : data <= 8'b00000000 ;
			12'h0000058E : data <= 8'b00000000 ;
			12'h0000058F : data <= 8'b00000000 ;
			12'h00000590 : data <= 8'b00000000 ;
			12'h00000591 : data <= 8'b00000000 ;
			12'h00000592 : data <= 8'b01100110 ;
			12'h00000593 : data <= 8'b01100110 ;
			12'h00000594 : data <= 8'b01100110 ;
			12'h00000595 : data <= 8'b01100110 ;
			12'h00000596 : data <= 8'b00111100 ;
			12'h00000597 : data <= 8'b00011000 ;
			12'h00000598 : data <= 8'b00011000 ;
			12'h00000599 : data <= 8'b00011000 ;
			12'h0000059A : data <= 8'b00011000 ;
			12'h0000059B : data <= 8'b00111100 ;
			12'h0000059C : data <= 8'b00000000 ;
			12'h0000059D : data <= 8'b00000000 ;
			12'h0000059E : data <= 8'b00000000 ;
			12'h0000059F : data <= 8'b00000000 ;
			12'h000005A0 : data <= 8'b00000000 ;
			12'h000005A1 : data <= 8'b00000000 ;
			12'h000005A2 : data <= 8'b11111110 ;
			12'h000005A3 : data <= 8'b11000110 ;
			12'h000005A4 : data <= 8'b10000110 ;
			12'h000005A5 : data <= 8'b00001100 ;
			12'h000005A6 : data <= 8'b00011000 ;
			12'h000005A7 : data <= 8'b00110000 ;
			12'h000005A8 : data <= 8'b01100000 ;
			12'h000005A9 : data <= 8'b11000010 ;
			12'h000005AA : data <= 8'b11000110 ;
			12'h000005AB : data <= 8'b11111110 ;
			12'h000005AC : data <= 8'b00000000 ;
			12'h000005AD : data <= 8'b00000000 ;
			12'h000005AE : data <= 8'b00000000 ;
			12'h000005AF : data <= 8'b00000000 ;
			12'h000005B0 : data <= 8'b00000000 ;
			12'h000005B1 : data <= 8'b00000000 ;
			12'h000005B2 : data <= 8'b00111100 ;
			12'h000005B3 : data <= 8'b00110000 ;
			12'h000005B4 : data <= 8'b00110000 ;
			12'h000005B5 : data <= 8'b00110000 ;
			12'h000005B6 : data <= 8'b00110000 ;
			12'h000005B7 : data <= 8'b00110000 ;
			12'h000005B8 : data <= 8'b00110000 ;
			12'h000005B9 : data <= 8'b00110000 ;
			12'h000005BA : data <= 8'b00110000 ;
			12'h000005BB : data <= 8'b00111100 ;
			12'h000005BC : data <= 8'b00000000 ;
			12'h000005BD : data <= 8'b00000000 ;
			12'h000005BE : data <= 8'b00000000 ;
			12'h000005BF : data <= 8'b00000000 ;
			12'h000005C0 : data <= 8'b00000000 ;
			12'h000005C1 : data <= 8'b00000000 ;
			12'h000005C2 : data <= 8'b00000000 ;
			12'h000005C3 : data <= 8'b10000000 ;
			12'h000005C4 : data <= 8'b11000000 ;
			12'h000005C5 : data <= 8'b11100000 ;
			12'h000005C6 : data <= 8'b01110000 ;
			12'h000005C7 : data <= 8'b00111000 ;
			12'h000005C8 : data <= 8'b00011100 ;
			12'h000005C9 : data <= 8'b00001110 ;
			12'h000005CA : data <= 8'b00000110 ;
			12'h000005CB : data <= 8'b00000010 ;
			12'h000005CC : data <= 8'b00000000 ;
			12'h000005CD : data <= 8'b00000000 ;
			12'h000005CE : data <= 8'b00000000 ;
			12'h000005CF : data <= 8'b00000000 ;
			12'h000005D0 : data <= 8'b00000000 ;
			12'h000005D1 : data <= 8'b00000000 ;
			12'h000005D2 : data <= 8'b00111100 ;
			12'h000005D3 : data <= 8'b00001100 ;
			12'h000005D4 : data <= 8'b00001100 ;
			12'h000005D5 : data <= 8'b00001100 ;
			12'h000005D6 : data <= 8'b00001100 ;
			12'h000005D7 : data <= 8'b00001100 ;
			12'h000005D8 : data <= 8'b00001100 ;
			12'h000005D9 : data <= 8'b00001100 ;
			12'h000005DA : data <= 8'b00001100 ;
			12'h000005DB : data <= 8'b00111100 ;
			12'h000005DC : data <= 8'b00000000 ;
			12'h000005DD : data <= 8'b00000000 ;
			12'h000005DE : data <= 8'b00000000 ;
			12'h000005DF : data <= 8'b00000000 ;
			12'h000005E0 : data <= 8'b00010000 ;
			12'h000005E1 : data <= 8'b00111000 ;
			12'h000005E2 : data <= 8'b01101100 ;
			12'h000005E3 : data <= 8'b11000110 ;
			12'h000005E4 : data <= 8'b00000000 ;
			12'h000005E5 : data <= 8'b00000000 ;
			12'h000005E6 : data <= 8'b00000000 ;
			12'h000005E7 : data <= 8'b00000000 ;
			12'h000005E8 : data <= 8'b00000000 ;
			12'h000005E9 : data <= 8'b00000000 ;
			12'h000005EA : data <= 8'b00000000 ;
			12'h000005EB : data <= 8'b00000000 ;
			12'h000005EC : data <= 8'b00000000 ;
			12'h000005ED : data <= 8'b00000000 ;
			12'h000005EE : data <= 8'b00000000 ;
			12'h000005EF : data <= 8'b00000000 ;
			12'h000005F0 : data <= 8'b00000000 ;
			12'h000005F1 : data <= 8'b00000000 ;
			12'h000005F2 : data <= 8'b00000000 ;
			12'h000005F3 : data <= 8'b00000000 ;
			12'h000005F4 : data <= 8'b00000000 ;
			12'h000005F5 : data <= 8'b00000000 ;
			12'h000005F6 : data <= 8'b00000000 ;
			12'h000005F7 : data <= 8'b00000000 ;
			12'h000005F8 : data <= 8'b00000000 ;
			12'h000005F9 : data <= 8'b00000000 ;
			12'h000005FA : data <= 8'b00000000 ;
			12'h000005FB : data <= 8'b00000000 ;
			12'h000005FC : data <= 8'b00000000 ;
			12'h000005FD : data <= 8'b11111111 ;
			12'h000005FE : data <= 8'b00000000 ;
			12'h000005FF : data <= 8'b00000000 ;
			12'h00000600 : data <= 8'b00110000 ;
			12'h00000601 : data <= 8'b00110000 ;
			12'h00000602 : data <= 8'b00011000 ;
			12'h00000603 : data <= 8'b00000000 ;
			12'h00000604 : data <= 8'b00000000 ;
			12'h00000605 : data <= 8'b00000000 ;
			12'h00000606 : data <= 8'b00000000 ;
			12'h00000607 : data <= 8'b00000000 ;
			12'h00000608 : data <= 8'b00000000 ;
			12'h00000609 : data <= 8'b00000000 ;
			12'h0000060A : data <= 8'b00000000 ;
			12'h0000060B : data <= 8'b00000000 ;
			12'h0000060C : data <= 8'b00000000 ;
			12'h0000060D : data <= 8'b00000000 ;
			12'h0000060E : data <= 8'b00000000 ;
			12'h0000060F : data <= 8'b00000000 ;
			12'h00000610 : data <= 8'b00000000 ;
			12'h00000611 : data <= 8'b00000000 ;
			12'h00000612 : data <= 8'b00000000 ;
			12'h00000613 : data <= 8'b00000000 ;
			12'h00000614 : data <= 8'b00000000 ;
			12'h00000615 : data <= 8'b01111000 ;
			12'h00000616 : data <= 8'b00001100 ;
			12'h00000617 : data <= 8'b01111100 ;
			12'h00000618 : data <= 8'b11001100 ;
			12'h00000619 : data <= 8'b11001100 ;
			12'h0000061A : data <= 8'b11001100 ;
			12'h0000061B : data <= 8'b01110110 ;
			12'h0000061C : data <= 8'b00000000 ;
			12'h0000061D : data <= 8'b00000000 ;
			12'h0000061E : data <= 8'b00000000 ;
			12'h0000061F : data <= 8'b00000000 ;
			12'h00000620 : data <= 8'b00000000 ;
			12'h00000621 : data <= 8'b00000000 ;
			12'h00000622 : data <= 8'b11100000 ;
			12'h00000623 : data <= 8'b01100000 ;
			12'h00000624 : data <= 8'b01100000 ;
			12'h00000625 : data <= 8'b01111000 ;
			12'h00000626 : data <= 8'b01101100 ;
			12'h00000627 : data <= 8'b01100110 ;
			12'h00000628 : data <= 8'b01100110 ;
			12'h00000629 : data <= 8'b01100110 ;
			12'h0000062A : data <= 8'b01100110 ;
			12'h0000062B : data <= 8'b01111100 ;
			12'h0000062C : data <= 8'b00000000 ;
			12'h0000062D : data <= 8'b00000000 ;
			12'h0000062E : data <= 8'b00000000 ;
			12'h0000062F : data <= 8'b00000000 ;
			12'h00000630 : data <= 8'b00000000 ;
			12'h00000631 : data <= 8'b00000000 ;
			12'h00000632 : data <= 8'b00000000 ;
			12'h00000633 : data <= 8'b00000000 ;
			12'h00000634 : data <= 8'b00000000 ;
			12'h00000635 : data <= 8'b01111100 ;
			12'h00000636 : data <= 8'b11000110 ;
			12'h00000637 : data <= 8'b11000000 ;
			12'h00000638 : data <= 8'b11000000 ;
			12'h00000639 : data <= 8'b11000000 ;
			12'h0000063A : data <= 8'b11000110 ;
			12'h0000063B : data <= 8'b01111100 ;
			12'h0000063C : data <= 8'b00000000 ;
			12'h0000063D : data <= 8'b00000000 ;
			12'h0000063E : data <= 8'b00000000 ;
			12'h0000063F : data <= 8'b00000000 ;
			12'h00000640 : data <= 8'b00000000 ;
			12'h00000641 : data <= 8'b00000000 ;
			12'h00000642 : data <= 8'b00011100 ;
			12'h00000643 : data <= 8'b00001100 ;
			12'h00000644 : data <= 8'b00001100 ;
			12'h00000645 : data <= 8'b00111100 ;
			12'h00000646 : data <= 8'b01101100 ;
			12'h00000647 : data <= 8'b11001100 ;
			12'h00000648 : data <= 8'b11001100 ;
			12'h00000649 : data <= 8'b11001100 ;
			12'h0000064A : data <= 8'b11001100 ;
			12'h0000064B : data <= 8'b01110110 ;
			12'h0000064C : data <= 8'b00000000 ;
			12'h0000064D : data <= 8'b00000000 ;
			12'h0000064E : data <= 8'b00000000 ;
			12'h0000064F : data <= 8'b00000000 ;
			12'h00000650 : data <= 8'b00000000 ;
			12'h00000651 : data <= 8'b00000000 ;
			12'h00000652 : data <= 8'b00000000 ;
			12'h00000653 : data <= 8'b00000000 ;
			12'h00000654 : data <= 8'b00000000 ;
			12'h00000655 : data <= 8'b01111100 ;
			12'h00000656 : data <= 8'b11000110 ;
			12'h00000657 : data <= 8'b11111110 ;
			12'h00000658 : data <= 8'b11000000 ;
			12'h00000659 : data <= 8'b11000000 ;
			12'h0000065A : data <= 8'b11000110 ;
			12'h0000065B : data <= 8'b01111100 ;
			12'h0000065C : data <= 8'b00000000 ;
			12'h0000065D : data <= 8'b00000000 ;
			12'h0000065E : data <= 8'b00000000 ;
			12'h0000065F : data <= 8'b00000000 ;
			12'h00000660 : data <= 8'b00000000 ;
			12'h00000661 : data <= 8'b00000000 ;
			12'h00000662 : data <= 8'b00111000 ;
			12'h00000663 : data <= 8'b01101100 ;
			12'h00000664 : data <= 8'b01100100 ;
			12'h00000665 : data <= 8'b01100000 ;
			12'h00000666 : data <= 8'b11110000 ;
			12'h00000667 : data <= 8'b01100000 ;
			12'h00000668 : data <= 8'b01100000 ;
			12'h00000669 : data <= 8'b01100000 ;
			12'h0000066A : data <= 8'b01100000 ;
			12'h0000066B : data <= 8'b11110000 ;
			12'h0000066C : data <= 8'b00000000 ;
			12'h0000066D : data <= 8'b00000000 ;
			12'h0000066E : data <= 8'b00000000 ;
			12'h0000066F : data <= 8'b00000000 ;
			12'h00000670 : data <= 8'b00000000 ;
			12'h00000671 : data <= 8'b00000000 ;
			12'h00000672 : data <= 8'b00000000 ;
			12'h00000673 : data <= 8'b00000000 ;
			12'h00000674 : data <= 8'b00000000 ;
			12'h00000675 : data <= 8'b01110110 ;
			12'h00000676 : data <= 8'b11001100 ;
			12'h00000677 : data <= 8'b11001100 ;
			12'h00000678 : data <= 8'b11001100 ;
			12'h00000679 : data <= 8'b11001100 ;
			12'h0000067A : data <= 8'b11001100 ;
			12'h0000067B : data <= 8'b01111100 ;
			12'h0000067C : data <= 8'b00001100 ;
			12'h0000067D : data <= 8'b11001100 ;
			12'h0000067E : data <= 8'b01111000 ;
			12'h0000067F : data <= 8'b00000000 ;
			12'h00000680 : data <= 8'b00000000 ;
			12'h00000681 : data <= 8'b00000000 ;
			12'h00000682 : data <= 8'b11100000 ;
			12'h00000683 : data <= 8'b01100000 ;
			12'h00000684 : data <= 8'b01100000 ;
			12'h00000685 : data <= 8'b01101100 ;
			12'h00000686 : data <= 8'b01110110 ;
			12'h00000687 : data <= 8'b01100110 ;
			12'h00000688 : data <= 8'b01100110 ;
			12'h00000689 : data <= 8'b01100110 ;
			12'h0000068A : data <= 8'b01100110 ;
			12'h0000068B : data <= 8'b11100110 ;
			12'h0000068C : data <= 8'b00000000 ;
			12'h0000068D : data <= 8'b00000000 ;
			12'h0000068E : data <= 8'b00000000 ;
			12'h0000068F : data <= 8'b00000000 ;
			12'h00000690 : data <= 8'b00000000 ;
			12'h00000691 : data <= 8'b00000000 ;
			12'h00000692 : data <= 8'b00011000 ;
			12'h00000693 : data <= 8'b00011000 ;
			12'h00000694 : data <= 8'b00000000 ;
			12'h00000695 : data <= 8'b00111000 ;
			12'h00000696 : data <= 8'b00011000 ;
			12'h00000697 : data <= 8'b00011000 ;
			12'h00000698 : data <= 8'b00011000 ;
			12'h00000699 : data <= 8'b00011000 ;
			12'h0000069A : data <= 8'b00011000 ;
			12'h0000069B : data <= 8'b00111100 ;
			12'h0000069C : data <= 8'b00000000 ;
			12'h0000069D : data <= 8'b00000000 ;
			12'h0000069E : data <= 8'b00000000 ;
			12'h0000069F : data <= 8'b00000000 ;
			12'h000006A0 : data <= 8'b00000000 ;
			12'h000006A1 : data <= 8'b00000000 ;
			12'h000006A2 : data <= 8'b00000110 ;
			12'h000006A3 : data <= 8'b00000110 ;
			12'h000006A4 : data <= 8'b00000000 ;
			12'h000006A5 : data <= 8'b00001110 ;
			12'h000006A6 : data <= 8'b00000110 ;
			12'h000006A7 : data <= 8'b00000110 ;
			12'h000006A8 : data <= 8'b00000110 ;
			12'h000006A9 : data <= 8'b00000110 ;
			12'h000006AA : data <= 8'b00000110 ;
			12'h000006AB : data <= 8'b00000110 ;
			12'h000006AC : data <= 8'b01100110 ;
			12'h000006AD : data <= 8'b01100110 ;
			12'h000006AE : data <= 8'b00111100 ;
			12'h000006AF : data <= 8'b00000000 ;
			12'h000006B0 : data <= 8'b00000000 ;
			12'h000006B1 : data <= 8'b00000000 ;
			12'h000006B2 : data <= 8'b11100000 ;
			12'h000006B3 : data <= 8'b01100000 ;
			12'h000006B4 : data <= 8'b01100000 ;
			12'h000006B5 : data <= 8'b01100110 ;
			12'h000006B6 : data <= 8'b01101100 ;
			12'h000006B7 : data <= 8'b01111000 ;
			12'h000006B8 : data <= 8'b01111000 ;
			12'h000006B9 : data <= 8'b01101100 ;
			12'h000006BA : data <= 8'b01100110 ;
			12'h000006BB : data <= 8'b11100110 ;
			12'h000006BC : data <= 8'b00000000 ;
			12'h000006BD : data <= 8'b00000000 ;
			12'h000006BE : data <= 8'b00000000 ;
			12'h000006BF : data <= 8'b00000000 ;
			12'h000006C0 : data <= 8'b00000000 ;
			12'h000006C1 : data <= 8'b00000000 ;
			12'h000006C2 : data <= 8'b00111000 ;
			12'h000006C3 : data <= 8'b00011000 ;
			12'h000006C4 : data <= 8'b00011000 ;
			12'h000006C5 : data <= 8'b00011000 ;
			12'h000006C6 : data <= 8'b00011000 ;
			12'h000006C7 : data <= 8'b00011000 ;
			12'h000006C8 : data <= 8'b00011000 ;
			12'h000006C9 : data <= 8'b00011000 ;
			12'h000006CA : data <= 8'b00011000 ;
			12'h000006CB : data <= 8'b00111100 ;
			12'h000006CC : data <= 8'b00000000 ;
			12'h000006CD : data <= 8'b00000000 ;
			12'h000006CE : data <= 8'b00000000 ;
			12'h000006CF : data <= 8'b00000000 ;
			12'h000006D0 : data <= 8'b00000000 ;
			12'h000006D1 : data <= 8'b00000000 ;
			12'h000006D2 : data <= 8'b00000000 ;
			12'h000006D3 : data <= 8'b00000000 ;
			12'h000006D4 : data <= 8'b00000000 ;
			12'h000006D5 : data <= 8'b11101100 ;
			12'h000006D6 : data <= 8'b11111110 ;
			12'h000006D7 : data <= 8'b11010110 ;
			12'h000006D8 : data <= 8'b11010110 ;
			12'h000006D9 : data <= 8'b11010110 ;
			12'h000006DA : data <= 8'b11010110 ;
			12'h000006DB : data <= 8'b11000110 ;
			12'h000006DC : data <= 8'b00000000 ;
			12'h000006DD : data <= 8'b00000000 ;
			12'h000006DE : data <= 8'b00000000 ;
			12'h000006DF : data <= 8'b00000000 ;
			12'h000006E0 : data <= 8'b00000000 ;
			12'h000006E1 : data <= 8'b00000000 ;
			12'h000006E2 : data <= 8'b00000000 ;
			12'h000006E3 : data <= 8'b00000000 ;
			12'h000006E4 : data <= 8'b00000000 ;
			12'h000006E5 : data <= 8'b11011100 ;
			12'h000006E6 : data <= 8'b01100110 ;
			12'h000006E7 : data <= 8'b01100110 ;
			12'h000006E8 : data <= 8'b01100110 ;
			12'h000006E9 : data <= 8'b01100110 ;
			12'h000006EA : data <= 8'b01100110 ;
			12'h000006EB : data <= 8'b01100110 ;
			12'h000006EC : data <= 8'b00000000 ;
			12'h000006ED : data <= 8'b00000000 ;
			12'h000006EE : data <= 8'b00000000 ;
			12'h000006EF : data <= 8'b00000000 ;
			12'h000006F0 : data <= 8'b00000000 ;
			12'h000006F1 : data <= 8'b00000000 ;
			12'h000006F2 : data <= 8'b00000000 ;
			12'h000006F3 : data <= 8'b00000000 ;
			12'h000006F4 : data <= 8'b00000000 ;
			12'h000006F5 : data <= 8'b01111100 ;
			12'h000006F6 : data <= 8'b11000110 ;
			12'h000006F7 : data <= 8'b11000110 ;
			12'h000006F8 : data <= 8'b11000110 ;
			12'h000006F9 : data <= 8'b11000110 ;
			12'h000006FA : data <= 8'b11000110 ;
			12'h000006FB : data <= 8'b01111100 ;
			12'h000006FC : data <= 8'b00000000 ;
			12'h000006FD : data <= 8'b00000000 ;
			12'h000006FE : data <= 8'b00000000 ;
			12'h000006FF : data <= 8'b00000000 ;
			12'h00000700 : data <= 8'b00000000 ;
			12'h00000701 : data <= 8'b00000000 ;
			12'h00000702 : data <= 8'b00000000 ;
			12'h00000703 : data <= 8'b00000000 ;
			12'h00000704 : data <= 8'b00000000 ;
			12'h00000705 : data <= 8'b11011100 ;
			12'h00000706 : data <= 8'b01100110 ;
			12'h00000707 : data <= 8'b01100110 ;
			12'h00000708 : data <= 8'b01100110 ;
			12'h00000709 : data <= 8'b01100110 ;
			12'h0000070A : data <= 8'b01100110 ;
			12'h0000070B : data <= 8'b01111100 ;
			12'h0000070C : data <= 8'b01100000 ;
			12'h0000070D : data <= 8'b01100000 ;
			12'h0000070E : data <= 8'b11110000 ;
			12'h0000070F : data <= 8'b00000000 ;
			12'h00000710 : data <= 8'b00000000 ;
			12'h00000711 : data <= 8'b00000000 ;
			12'h00000712 : data <= 8'b00000000 ;
			12'h00000713 : data <= 8'b00000000 ;
			12'h00000714 : data <= 8'b00000000 ;
			12'h00000715 : data <= 8'b01110110 ;
			12'h00000716 : data <= 8'b11001100 ;
			12'h00000717 : data <= 8'b11001100 ;
			12'h00000718 : data <= 8'b11001100 ;
			12'h00000719 : data <= 8'b11001100 ;
			12'h0000071A : data <= 8'b11001100 ;
			12'h0000071B : data <= 8'b01111100 ;
			12'h0000071C : data <= 8'b00001100 ;
			12'h0000071D : data <= 8'b00001100 ;
			12'h0000071E : data <= 8'b00011110 ;
			12'h0000071F : data <= 8'b00000000 ;
			12'h00000720 : data <= 8'b00000000 ;
			12'h00000721 : data <= 8'b00000000 ;
			12'h00000722 : data <= 8'b00000000 ;
			12'h00000723 : data <= 8'b00000000 ;
			12'h00000724 : data <= 8'b00000000 ;
			12'h00000725 : data <= 8'b11011100 ;
			12'h00000726 : data <= 8'b01110110 ;
			12'h00000727 : data <= 8'b01100110 ;
			12'h00000728 : data <= 8'b01100000 ;
			12'h00000729 : data <= 8'b01100000 ;
			12'h0000072A : data <= 8'b01100000 ;
			12'h0000072B : data <= 8'b11110000 ;
			12'h0000072C : data <= 8'b00000000 ;
			12'h0000072D : data <= 8'b00000000 ;
			12'h0000072E : data <= 8'b00000000 ;
			12'h0000072F : data <= 8'b00000000 ;
			12'h00000730 : data <= 8'b00000000 ;
			12'h00000731 : data <= 8'b00000000 ;
			12'h00000732 : data <= 8'b00000000 ;
			12'h00000733 : data <= 8'b00000000 ;
			12'h00000734 : data <= 8'b00000000 ;
			12'h00000735 : data <= 8'b01111100 ;
			12'h00000736 : data <= 8'b11000110 ;
			12'h00000737 : data <= 8'b01100000 ;
			12'h00000738 : data <= 8'b00111000 ;
			12'h00000739 : data <= 8'b00001100 ;
			12'h0000073A : data <= 8'b11000110 ;
			12'h0000073B : data <= 8'b01111100 ;
			12'h0000073C : data <= 8'b00000000 ;
			12'h0000073D : data <= 8'b00000000 ;
			12'h0000073E : data <= 8'b00000000 ;
			12'h0000073F : data <= 8'b00000000 ;
			12'h00000740 : data <= 8'b00000000 ;
			12'h00000741 : data <= 8'b00000000 ;
			12'h00000742 : data <= 8'b00010000 ;
			12'h00000743 : data <= 8'b00110000 ;
			12'h00000744 : data <= 8'b00110000 ;
			12'h00000745 : data <= 8'b11111100 ;
			12'h00000746 : data <= 8'b00110000 ;
			12'h00000747 : data <= 8'b00110000 ;
			12'h00000748 : data <= 8'b00110000 ;
			12'h00000749 : data <= 8'b00110000 ;
			12'h0000074A : data <= 8'b00110110 ;
			12'h0000074B : data <= 8'b00011100 ;
			12'h0000074C : data <= 8'b00000000 ;
			12'h0000074D : data <= 8'b00000000 ;
			12'h0000074E : data <= 8'b00000000 ;
			12'h0000074F : data <= 8'b00000000 ;
			12'h00000750 : data <= 8'b00000000 ;
			12'h00000751 : data <= 8'b00000000 ;
			12'h00000752 : data <= 8'b00000000 ;
			12'h00000753 : data <= 8'b00000000 ;
			12'h00000754 : data <= 8'b00000000 ;
			12'h00000755 : data <= 8'b11001100 ;
			12'h00000756 : data <= 8'b11001100 ;
			12'h00000757 : data <= 8'b11001100 ;
			12'h00000758 : data <= 8'b11001100 ;
			12'h00000759 : data <= 8'b11001100 ;
			12'h0000075A : data <= 8'b11001100 ;
			12'h0000075B : data <= 8'b01110110 ;
			12'h0000075C : data <= 8'b00000000 ;
			12'h0000075D : data <= 8'b00000000 ;
			12'h0000075E : data <= 8'b00000000 ;
			12'h0000075F : data <= 8'b00000000 ;
			12'h00000760 : data <= 8'b00000000 ;
			12'h00000761 : data <= 8'b00000000 ;
			12'h00000762 : data <= 8'b00000000 ;
			12'h00000763 : data <= 8'b00000000 ;
			12'h00000764 : data <= 8'b00000000 ;
			12'h00000765 : data <= 8'b01100110 ;
			12'h00000766 : data <= 8'b01100110 ;
			12'h00000767 : data <= 8'b01100110 ;
			12'h00000768 : data <= 8'b01100110 ;
			12'h00000769 : data <= 8'b01100110 ;
			12'h0000076A : data <= 8'b00111100 ;
			12'h0000076B : data <= 8'b00011000 ;
			12'h0000076C : data <= 8'b00000000 ;
			12'h0000076D : data <= 8'b00000000 ;
			12'h0000076E : data <= 8'b00000000 ;
			12'h0000076F : data <= 8'b00000000 ;
			12'h00000770 : data <= 8'b00000000 ;
			12'h00000771 : data <= 8'b00000000 ;
			12'h00000772 : data <= 8'b00000000 ;
			12'h00000773 : data <= 8'b00000000 ;
			12'h00000774 : data <= 8'b00000000 ;
			12'h00000775 : data <= 8'b11000110 ;
			12'h00000776 : data <= 8'b11000110 ;
			12'h00000777 : data <= 8'b11010110 ;
			12'h00000778 : data <= 8'b11010110 ;
			12'h00000779 : data <= 8'b11010110 ;
			12'h0000077A : data <= 8'b11111110 ;
			12'h0000077B : data <= 8'b01101100 ;
			12'h0000077C : data <= 8'b00000000 ;
			12'h0000077D : data <= 8'b00000000 ;
			12'h0000077E : data <= 8'b00000000 ;
			12'h0000077F : data <= 8'b00000000 ;
			12'h00000780 : data <= 8'b00000000 ;
			12'h00000781 : data <= 8'b00000000 ;
			12'h00000782 : data <= 8'b00000000 ;
			12'h00000783 : data <= 8'b00000000 ;
			12'h00000784 : data <= 8'b00000000 ;
			12'h00000785 : data <= 8'b11000110 ;
			12'h00000786 : data <= 8'b01101100 ;
			12'h00000787 : data <= 8'b00111000 ;
			12'h00000788 : data <= 8'b00111000 ;
			12'h00000789 : data <= 8'b00111000 ;
			12'h0000078A : data <= 8'b01101100 ;
			12'h0000078B : data <= 8'b11000110 ;
			12'h0000078C : data <= 8'b00000000 ;
			12'h0000078D : data <= 8'b00000000 ;
			12'h0000078E : data <= 8'b00000000 ;
			12'h0000078F : data <= 8'b00000000 ;
			12'h00000790 : data <= 8'b00000000 ;
			12'h00000791 : data <= 8'b00000000 ;
			12'h00000792 : data <= 8'b00000000 ;
			12'h00000793 : data <= 8'b00000000 ;
			12'h00000794 : data <= 8'b00000000 ;
			12'h00000795 : data <= 8'b11000110 ;
			12'h00000796 : data <= 8'b11000110 ;
			12'h00000797 : data <= 8'b11000110 ;
			12'h00000798 : data <= 8'b11000110 ;
			12'h00000799 : data <= 8'b11000110 ;
			12'h0000079A : data <= 8'b11000110 ;
			12'h0000079B : data <= 8'b01111110 ;
			12'h0000079C : data <= 8'b00000110 ;
			12'h0000079D : data <= 8'b00001100 ;
			12'h0000079E : data <= 8'b11111000 ;
			12'h0000079F : data <= 8'b00000000 ;
			12'h000007A0 : data <= 8'b00000000 ;
			12'h000007A1 : data <= 8'b00000000 ;
			12'h000007A2 : data <= 8'b00000000 ;
			12'h000007A3 : data <= 8'b00000000 ;
			12'h000007A4 : data <= 8'b00000000 ;
			12'h000007A5 : data <= 8'b11111110 ;
			12'h000007A6 : data <= 8'b11001100 ;
			12'h000007A7 : data <= 8'b00011000 ;
			12'h000007A8 : data <= 8'b00110000 ;
			12'h000007A9 : data <= 8'b01100000 ;
			12'h000007AA : data <= 8'b11000110 ;
			12'h000007AB : data <= 8'b11111110 ;
			12'h000007AC : data <= 8'b00000000 ;
			12'h000007AD : data <= 8'b00000000 ;
			12'h000007AE : data <= 8'b00000000 ;
			12'h000007AF : data <= 8'b00000000 ;
			12'h000007B0 : data <= 8'b00000000 ;
			12'h000007B1 : data <= 8'b00000000 ;
			12'h000007B2 : data <= 8'b00001110 ;
			12'h000007B3 : data <= 8'b00011000 ;
			12'h000007B4 : data <= 8'b00011000 ;
			12'h000007B5 : data <= 8'b00011000 ;
			12'h000007B6 : data <= 8'b01110000 ;
			12'h000007B7 : data <= 8'b00011000 ;
			12'h000007B8 : data <= 8'b00011000 ;
			12'h000007B9 : data <= 8'b00011000 ;
			12'h000007BA : data <= 8'b00011000 ;
			12'h000007BB : data <= 8'b00001110 ;
			12'h000007BC : data <= 8'b00000000 ;
			12'h000007BD : data <= 8'b00000000 ;
			12'h000007BE : data <= 8'b00000000 ;
			12'h000007BF : data <= 8'b00000000 ;
			12'h000007C0 : data <= 8'b00000000 ;
			12'h000007C1 : data <= 8'b00000000 ;
			12'h000007C2 : data <= 8'b00011000 ;
			12'h000007C3 : data <= 8'b00011000 ;
			12'h000007C4 : data <= 8'b00011000 ;
			12'h000007C5 : data <= 8'b00011000 ;
			12'h000007C6 : data <= 8'b00000000 ;
			12'h000007C7 : data <= 8'b00011000 ;
			12'h000007C8 : data <= 8'b00011000 ;
			12'h000007C9 : data <= 8'b00011000 ;
			12'h000007CA : data <= 8'b00011000 ;
			12'h000007CB : data <= 8'b00011000 ;
			12'h000007CC : data <= 8'b00000000 ;
			12'h000007CD : data <= 8'b00000000 ;
			12'h000007CE : data <= 8'b00000000 ;
			12'h000007CF : data <= 8'b00000000 ;
			12'h000007D0 : data <= 8'b00000000 ;
			12'h000007D1 : data <= 8'b00000000 ;
			12'h000007D2 : data <= 8'b01110000 ;
			12'h000007D3 : data <= 8'b00011000 ;
			12'h000007D4 : data <= 8'b00011000 ;
			12'h000007D5 : data <= 8'b00011000 ;
			12'h000007D6 : data <= 8'b00001110 ;
			12'h000007D7 : data <= 8'b00011000 ;
			12'h000007D8 : data <= 8'b00011000 ;
			12'h000007D9 : data <= 8'b00011000 ;
			12'h000007DA : data <= 8'b00011000 ;
			12'h000007DB : data <= 8'b01110000 ;
			12'h000007DC : data <= 8'b00000000 ;
			12'h000007DD : data <= 8'b00000000 ;
			12'h000007DE : data <= 8'b00000000 ;
			12'h000007DF : data <= 8'b00000000 ;
			12'h000007E0 : data <= 8'b00000000 ;
			12'h000007E1 : data <= 8'b00000000 ;
			12'h000007E2 : data <= 8'b01110110 ;
			12'h000007E3 : data <= 8'b11011100 ;
			12'h000007E4 : data <= 8'b00000000 ;
			12'h000007E5 : data <= 8'b00000000 ;
			12'h000007E6 : data <= 8'b00000000 ;
			12'h000007E7 : data <= 8'b00000000 ;
			12'h000007E8 : data <= 8'b00000000 ;
			12'h000007E9 : data <= 8'b00000000 ;
			12'h000007EA : data <= 8'b00000000 ;
			12'h000007EB : data <= 8'b00000000 ;
			12'h000007EC : data <= 8'b00000000 ;
			12'h000007ED : data <= 8'b00000000 ;
			12'h000007EE : data <= 8'b00000000 ;
			12'h000007EF : data <= 8'b00000000 ;
			12'h000007F0 : data <= 8'b00000000 ;
			12'h000007F1 : data <= 8'b00000000 ;
			12'h000007F2 : data <= 8'b00000000 ;
			12'h000007F3 : data <= 8'b00000000 ;
			12'h000007F4 : data <= 8'b00010000 ;
			12'h000007F5 : data <= 8'b00111000 ;
			12'h000007F6 : data <= 8'b01101100 ;
			12'h000007F7 : data <= 8'b11000110 ;
			12'h000007F8 : data <= 8'b11000110 ;
			12'h000007F9 : data <= 8'b11000110 ;
			12'h000007FA : data <= 8'b11111110 ;
			12'h000007FB : data <= 8'b00000000 ;
			12'h000007FC : data <= 8'b00000000 ;
			12'h000007FD : data <= 8'b00000000 ;
			12'h000007FE : data <= 8'b00000000 ;
			12'h000007FF : data <= 8'b00000000 ;
			12'h00000800 : data <= 8'b00000000 ;
			12'h00000801 : data <= 8'b00000000 ;
			12'h00000802 : data <= 8'b00111100 ;
			12'h00000803 : data <= 8'b01100110 ;
			12'h00000804 : data <= 8'b11000010 ;
			12'h00000805 : data <= 8'b11000000 ;
			12'h00000806 : data <= 8'b11000000 ;
			12'h00000807 : data <= 8'b11000000 ;
			12'h00000808 : data <= 8'b11000010 ;
			12'h00000809 : data <= 8'b01100110 ;
			12'h0000080A : data <= 8'b00111100 ;
			12'h0000080B : data <= 8'b00001100 ;
			12'h0000080C : data <= 8'b00000110 ;
			12'h0000080D : data <= 8'b01111100 ;
			12'h0000080E : data <= 8'b00000000 ;
			12'h0000080F : data <= 8'b00000000 ;
			12'h00000810 : data <= 8'b00000000 ;
			12'h00000811 : data <= 8'b00000000 ;
			12'h00000812 : data <= 8'b11001100 ;
			12'h00000813 : data <= 8'b00000000 ;
			12'h00000814 : data <= 8'b00000000 ;
			12'h00000815 : data <= 8'b11001100 ;
			12'h00000816 : data <= 8'b11001100 ;
			12'h00000817 : data <= 8'b11001100 ;
			12'h00000818 : data <= 8'b11001100 ;
			12'h00000819 : data <= 8'b11001100 ;
			12'h0000081A : data <= 8'b11001100 ;
			12'h0000081B : data <= 8'b01110110 ;
			12'h0000081C : data <= 8'b00000000 ;
			12'h0000081D : data <= 8'b00000000 ;
			12'h0000081E : data <= 8'b00000000 ;
			12'h0000081F : data <= 8'b00000000 ;
			12'h00000820 : data <= 8'b00000000 ;
			12'h00000821 : data <= 8'b00001100 ;
			12'h00000822 : data <= 8'b00011000 ;
			12'h00000823 : data <= 8'b00110000 ;
			12'h00000824 : data <= 8'b00000000 ;
			12'h00000825 : data <= 8'b01111100 ;
			12'h00000826 : data <= 8'b11000110 ;
			12'h00000827 : data <= 8'b11111110 ;
			12'h00000828 : data <= 8'b11000000 ;
			12'h00000829 : data <= 8'b11000000 ;
			12'h0000082A : data <= 8'b11000110 ;
			12'h0000082B : data <= 8'b01111100 ;
			12'h0000082C : data <= 8'b00000000 ;
			12'h0000082D : data <= 8'b00000000 ;
			12'h0000082E : data <= 8'b00000000 ;
			12'h0000082F : data <= 8'b00000000 ;
			12'h00000830 : data <= 8'b00000000 ;
			12'h00000831 : data <= 8'b00010000 ;
			12'h00000832 : data <= 8'b00111000 ;
			12'h00000833 : data <= 8'b01101100 ;
			12'h00000834 : data <= 8'b00000000 ;
			12'h00000835 : data <= 8'b01111000 ;
			12'h00000836 : data <= 8'b00001100 ;
			12'h00000837 : data <= 8'b01111100 ;
			12'h00000838 : data <= 8'b11001100 ;
			12'h00000839 : data <= 8'b11001100 ;
			12'h0000083A : data <= 8'b11001100 ;
			12'h0000083B : data <= 8'b01110110 ;
			12'h0000083C : data <= 8'b00000000 ;
			12'h0000083D : data <= 8'b00000000 ;
			12'h0000083E : data <= 8'b00000000 ;
			12'h0000083F : data <= 8'b00000000 ;
			12'h00000840 : data <= 8'b00000000 ;
			12'h00000841 : data <= 8'b00000000 ;
			12'h00000842 : data <= 8'b11001100 ;
			12'h00000843 : data <= 8'b00000000 ;
			12'h00000844 : data <= 8'b00000000 ;
			12'h00000845 : data <= 8'b01111000 ;
			12'h00000846 : data <= 8'b00001100 ;
			12'h00000847 : data <= 8'b01111100 ;
			12'h00000848 : data <= 8'b11001100 ;
			12'h00000849 : data <= 8'b11001100 ;
			12'h0000084A : data <= 8'b11001100 ;
			12'h0000084B : data <= 8'b01110110 ;
			12'h0000084C : data <= 8'b00000000 ;
			12'h0000084D : data <= 8'b00000000 ;
			12'h0000084E : data <= 8'b00000000 ;
			12'h0000084F : data <= 8'b00000000 ;
			12'h00000850 : data <= 8'b00000000 ;
			12'h00000851 : data <= 8'b01100000 ;
			12'h00000852 : data <= 8'b00110000 ;
			12'h00000853 : data <= 8'b00011000 ;
			12'h00000854 : data <= 8'b00000000 ;
			12'h00000855 : data <= 8'b01111000 ;
			12'h00000856 : data <= 8'b00001100 ;
			12'h00000857 : data <= 8'b01111100 ;
			12'h00000858 : data <= 8'b11001100 ;
			12'h00000859 : data <= 8'b11001100 ;
			12'h0000085A : data <= 8'b11001100 ;
			12'h0000085B : data <= 8'b01110110 ;
			12'h0000085C : data <= 8'b00000000 ;
			12'h0000085D : data <= 8'b00000000 ;
			12'h0000085E : data <= 8'b00000000 ;
			12'h0000085F : data <= 8'b00000000 ;
			12'h00000860 : data <= 8'b00000000 ;
			12'h00000861 : data <= 8'b00111000 ;
			12'h00000862 : data <= 8'b01101100 ;
			12'h00000863 : data <= 8'b00111000 ;
			12'h00000864 : data <= 8'b00000000 ;
			12'h00000865 : data <= 8'b01111000 ;
			12'h00000866 : data <= 8'b00001100 ;
			12'h00000867 : data <= 8'b01111100 ;
			12'h00000868 : data <= 8'b11001100 ;
			12'h00000869 : data <= 8'b11001100 ;
			12'h0000086A : data <= 8'b11001100 ;
			12'h0000086B : data <= 8'b01110110 ;
			12'h0000086C : data <= 8'b00000000 ;
			12'h0000086D : data <= 8'b00000000 ;
			12'h0000086E : data <= 8'b00000000 ;
			12'h0000086F : data <= 8'b00000000 ;
			12'h00000870 : data <= 8'b00000000 ;
			12'h00000871 : data <= 8'b00000000 ;
			12'h00000872 : data <= 8'b00000000 ;
			12'h00000873 : data <= 8'b00000000 ;
			12'h00000874 : data <= 8'b00111100 ;
			12'h00000875 : data <= 8'b01100110 ;
			12'h00000876 : data <= 8'b01100000 ;
			12'h00000877 : data <= 8'b01100000 ;
			12'h00000878 : data <= 8'b01100110 ;
			12'h00000879 : data <= 8'b00111100 ;
			12'h0000087A : data <= 8'b00001100 ;
			12'h0000087B : data <= 8'b00000110 ;
			12'h0000087C : data <= 8'b00111100 ;
			12'h0000087D : data <= 8'b00000000 ;
			12'h0000087E : data <= 8'b00000000 ;
			12'h0000087F : data <= 8'b00000000 ;
			12'h00000880 : data <= 8'b00000000 ;
			12'h00000881 : data <= 8'b00010000 ;
			12'h00000882 : data <= 8'b00111000 ;
			12'h00000883 : data <= 8'b01101100 ;
			12'h00000884 : data <= 8'b00000000 ;
			12'h00000885 : data <= 8'b01111100 ;
			12'h00000886 : data <= 8'b11000110 ;
			12'h00000887 : data <= 8'b11111110 ;
			12'h00000888 : data <= 8'b11000000 ;
			12'h00000889 : data <= 8'b11000000 ;
			12'h0000088A : data <= 8'b11000110 ;
			12'h0000088B : data <= 8'b01111100 ;
			12'h0000088C : data <= 8'b00000000 ;
			12'h0000088D : data <= 8'b00000000 ;
			12'h0000088E : data <= 8'b00000000 ;
			12'h0000088F : data <= 8'b00000000 ;
			12'h00000890 : data <= 8'b00000000 ;
			12'h00000891 : data <= 8'b00000000 ;
			12'h00000892 : data <= 8'b11000110 ;
			12'h00000893 : data <= 8'b00000000 ;
			12'h00000894 : data <= 8'b00000000 ;
			12'h00000895 : data <= 8'b01111100 ;
			12'h00000896 : data <= 8'b11000110 ;
			12'h00000897 : data <= 8'b11111110 ;
			12'h00000898 : data <= 8'b11000000 ;
			12'h00000899 : data <= 8'b11000000 ;
			12'h0000089A : data <= 8'b11000110 ;
			12'h0000089B : data <= 8'b01111100 ;
			12'h0000089C : data <= 8'b00000000 ;
			12'h0000089D : data <= 8'b00000000 ;
			12'h0000089E : data <= 8'b00000000 ;
			12'h0000089F : data <= 8'b00000000 ;
			12'h000008A0 : data <= 8'b00000000 ;
			12'h000008A1 : data <= 8'b01100000 ;
			12'h000008A2 : data <= 8'b00110000 ;
			12'h000008A3 : data <= 8'b00011000 ;
			12'h000008A4 : data <= 8'b00000000 ;
			12'h000008A5 : data <= 8'b01111100 ;
			12'h000008A6 : data <= 8'b11000110 ;
			12'h000008A7 : data <= 8'b11111110 ;
			12'h000008A8 : data <= 8'b11000000 ;
			12'h000008A9 : data <= 8'b11000000 ;
			12'h000008AA : data <= 8'b11000110 ;
			12'h000008AB : data <= 8'b01111100 ;
			12'h000008AC : data <= 8'b00000000 ;
			12'h000008AD : data <= 8'b00000000 ;
			12'h000008AE : data <= 8'b00000000 ;
			12'h000008AF : data <= 8'b00000000 ;
			12'h000008B0 : data <= 8'b00000000 ;
			12'h000008B1 : data <= 8'b00000000 ;
			12'h000008B2 : data <= 8'b01100110 ;
			12'h000008B3 : data <= 8'b00000000 ;
			12'h000008B4 : data <= 8'b00000000 ;
			12'h000008B5 : data <= 8'b00111000 ;
			12'h000008B6 : data <= 8'b00011000 ;
			12'h000008B7 : data <= 8'b00011000 ;
			12'h000008B8 : data <= 8'b00011000 ;
			12'h000008B9 : data <= 8'b00011000 ;
			12'h000008BA : data <= 8'b00011000 ;
			12'h000008BB : data <= 8'b00111100 ;
			12'h000008BC : data <= 8'b00000000 ;
			12'h000008BD : data <= 8'b00000000 ;
			12'h000008BE : data <= 8'b00000000 ;
			12'h000008BF : data <= 8'b00000000 ;
			12'h000008C0 : data <= 8'b00000000 ;
			12'h000008C1 : data <= 8'b00011000 ;
			12'h000008C2 : data <= 8'b00111100 ;
			12'h000008C3 : data <= 8'b01100110 ;
			12'h000008C4 : data <= 8'b00000000 ;
			12'h000008C5 : data <= 8'b00111000 ;
			12'h000008C6 : data <= 8'b00011000 ;
			12'h000008C7 : data <= 8'b00011000 ;
			12'h000008C8 : data <= 8'b00011000 ;
			12'h000008C9 : data <= 8'b00011000 ;
			12'h000008CA : data <= 8'b00011000 ;
			12'h000008CB : data <= 8'b00111100 ;
			12'h000008CC : data <= 8'b00000000 ;
			12'h000008CD : data <= 8'b00000000 ;
			12'h000008CE : data <= 8'b00000000 ;
			12'h000008CF : data <= 8'b00000000 ;
			12'h000008D0 : data <= 8'b00000000 ;
			12'h000008D1 : data <= 8'b01100000 ;
			12'h000008D2 : data <= 8'b00110000 ;
			12'h000008D3 : data <= 8'b00011000 ;
			12'h000008D4 : data <= 8'b00000000 ;
			12'h000008D5 : data <= 8'b00111000 ;
			12'h000008D6 : data <= 8'b00011000 ;
			12'h000008D7 : data <= 8'b00011000 ;
			12'h000008D8 : data <= 8'b00011000 ;
			12'h000008D9 : data <= 8'b00011000 ;
			12'h000008DA : data <= 8'b00011000 ;
			12'h000008DB : data <= 8'b00111100 ;
			12'h000008DC : data <= 8'b00000000 ;
			12'h000008DD : data <= 8'b00000000 ;
			12'h000008DE : data <= 8'b00000000 ;
			12'h000008DF : data <= 8'b00000000 ;
			12'h000008E0 : data <= 8'b00000000 ;
			12'h000008E1 : data <= 8'b11000110 ;
			12'h000008E2 : data <= 8'b00000000 ;
			12'h000008E3 : data <= 8'b00010000 ;
			12'h000008E4 : data <= 8'b00111000 ;
			12'h000008E5 : data <= 8'b01101100 ;
			12'h000008E6 : data <= 8'b11000110 ;
			12'h000008E7 : data <= 8'b11000110 ;
			12'h000008E8 : data <= 8'b11111110 ;
			12'h000008E9 : data <= 8'b11000110 ;
			12'h000008EA : data <= 8'b11000110 ;
			12'h000008EB : data <= 8'b11000110 ;
			12'h000008EC : data <= 8'b00000000 ;
			12'h000008ED : data <= 8'b00000000 ;
			12'h000008EE : data <= 8'b00000000 ;
			12'h000008EF : data <= 8'b00000000 ;
			12'h000008F0 : data <= 8'b00111000 ;
			12'h000008F1 : data <= 8'b01101100 ;
			12'h000008F2 : data <= 8'b00111000 ;
			12'h000008F3 : data <= 8'b00000000 ;
			12'h000008F4 : data <= 8'b00111000 ;
			12'h000008F5 : data <= 8'b01101100 ;
			12'h000008F6 : data <= 8'b11000110 ;
			12'h000008F7 : data <= 8'b11000110 ;
			12'h000008F8 : data <= 8'b11111110 ;
			12'h000008F9 : data <= 8'b11000110 ;
			12'h000008FA : data <= 8'b11000110 ;
			12'h000008FB : data <= 8'b11000110 ;
			12'h000008FC : data <= 8'b00000000 ;
			12'h000008FD : data <= 8'b00000000 ;
			12'h000008FE : data <= 8'b00000000 ;
			12'h000008FF : data <= 8'b00000000 ;
			12'h00000900 : data <= 8'b00011000 ;
			12'h00000901 : data <= 8'b00110000 ;
			12'h00000902 : data <= 8'b01100000 ;
			12'h00000903 : data <= 8'b00000000 ;
			12'h00000904 : data <= 8'b11111110 ;
			12'h00000905 : data <= 8'b01100110 ;
			12'h00000906 : data <= 8'b01100000 ;
			12'h00000907 : data <= 8'b01111100 ;
			12'h00000908 : data <= 8'b01100000 ;
			12'h00000909 : data <= 8'b01100000 ;
			12'h0000090A : data <= 8'b01100110 ;
			12'h0000090B : data <= 8'b11111110 ;
			12'h0000090C : data <= 8'b00000000 ;
			12'h0000090D : data <= 8'b00000000 ;
			12'h0000090E : data <= 8'b00000000 ;
			12'h0000090F : data <= 8'b00000000 ;
			12'h00000910 : data <= 8'b00000000 ;
			12'h00000911 : data <= 8'b00000000 ;
			12'h00000912 : data <= 8'b00000000 ;
			12'h00000913 : data <= 8'b00000000 ;
			12'h00000914 : data <= 8'b00000000 ;
			12'h00000915 : data <= 8'b11001100 ;
			12'h00000916 : data <= 8'b01110110 ;
			12'h00000917 : data <= 8'b00110110 ;
			12'h00000918 : data <= 8'b01111110 ;
			12'h00000919 : data <= 8'b11011000 ;
			12'h0000091A : data <= 8'b11011000 ;
			12'h0000091B : data <= 8'b01101110 ;
			12'h0000091C : data <= 8'b00000000 ;
			12'h0000091D : data <= 8'b00000000 ;
			12'h0000091E : data <= 8'b00000000 ;
			12'h0000091F : data <= 8'b00000000 ;
			12'h00000920 : data <= 8'b00000000 ;
			12'h00000921 : data <= 8'b00000000 ;
			12'h00000922 : data <= 8'b00111110 ;
			12'h00000923 : data <= 8'b01101100 ;
			12'h00000924 : data <= 8'b11001100 ;
			12'h00000925 : data <= 8'b11001100 ;
			12'h00000926 : data <= 8'b11111110 ;
			12'h00000927 : data <= 8'b11001100 ;
			12'h00000928 : data <= 8'b11001100 ;
			12'h00000929 : data <= 8'b11001100 ;
			12'h0000092A : data <= 8'b11001100 ;
			12'h0000092B : data <= 8'b11001110 ;
			12'h0000092C : data <= 8'b00000000 ;
			12'h0000092D : data <= 8'b00000000 ;
			12'h0000092E : data <= 8'b00000000 ;
			12'h0000092F : data <= 8'b00000000 ;
			12'h00000930 : data <= 8'b00000000 ;
			12'h00000931 : data <= 8'b00010000 ;
			12'h00000932 : data <= 8'b00111000 ;
			12'h00000933 : data <= 8'b01101100 ;
			12'h00000934 : data <= 8'b00000000 ;
			12'h00000935 : data <= 8'b01111100 ;
			12'h00000936 : data <= 8'b11000110 ;
			12'h00000937 : data <= 8'b11000110 ;
			12'h00000938 : data <= 8'b11000110 ;
			12'h00000939 : data <= 8'b11000110 ;
			12'h0000093A : data <= 8'b11000110 ;
			12'h0000093B : data <= 8'b01111100 ;
			12'h0000093C : data <= 8'b00000000 ;
			12'h0000093D : data <= 8'b00000000 ;
			12'h0000093E : data <= 8'b00000000 ;
			12'h0000093F : data <= 8'b00000000 ;
			12'h00000940 : data <= 8'b00000000 ;
			12'h00000941 : data <= 8'b00000000 ;
			12'h00000942 : data <= 8'b11000110 ;
			12'h00000943 : data <= 8'b00000000 ;
			12'h00000944 : data <= 8'b00000000 ;
			12'h00000945 : data <= 8'b01111100 ;
			12'h00000946 : data <= 8'b11000110 ;
			12'h00000947 : data <= 8'b11000110 ;
			12'h00000948 : data <= 8'b11000110 ;
			12'h00000949 : data <= 8'b11000110 ;
			12'h0000094A : data <= 8'b11000110 ;
			12'h0000094B : data <= 8'b01111100 ;
			12'h0000094C : data <= 8'b00000000 ;
			12'h0000094D : data <= 8'b00000000 ;
			12'h0000094E : data <= 8'b00000000 ;
			12'h0000094F : data <= 8'b00000000 ;
			12'h00000950 : data <= 8'b00000000 ;
			12'h00000951 : data <= 8'b01100000 ;
			12'h00000952 : data <= 8'b00110000 ;
			12'h00000953 : data <= 8'b00011000 ;
			12'h00000954 : data <= 8'b00000000 ;
			12'h00000955 : data <= 8'b01111100 ;
			12'h00000956 : data <= 8'b11000110 ;
			12'h00000957 : data <= 8'b11000110 ;
			12'h00000958 : data <= 8'b11000110 ;
			12'h00000959 : data <= 8'b11000110 ;
			12'h0000095A : data <= 8'b11000110 ;
			12'h0000095B : data <= 8'b01111100 ;
			12'h0000095C : data <= 8'b00000000 ;
			12'h0000095D : data <= 8'b00000000 ;
			12'h0000095E : data <= 8'b00000000 ;
			12'h0000095F : data <= 8'b00000000 ;
			12'h00000960 : data <= 8'b00000000 ;
			12'h00000961 : data <= 8'b00110000 ;
			12'h00000962 : data <= 8'b01111000 ;
			12'h00000963 : data <= 8'b11001100 ;
			12'h00000964 : data <= 8'b00000000 ;
			12'h00000965 : data <= 8'b11001100 ;
			12'h00000966 : data <= 8'b11001100 ;
			12'h00000967 : data <= 8'b11001100 ;
			12'h00000968 : data <= 8'b11001100 ;
			12'h00000969 : data <= 8'b11001100 ;
			12'h0000096A : data <= 8'b11001100 ;
			12'h0000096B : data <= 8'b01110110 ;
			12'h0000096C : data <= 8'b00000000 ;
			12'h0000096D : data <= 8'b00000000 ;
			12'h0000096E : data <= 8'b00000000 ;
			12'h0000096F : data <= 8'b00000000 ;
			12'h00000970 : data <= 8'b00000000 ;
			12'h00000971 : data <= 8'b01100000 ;
			12'h00000972 : data <= 8'b00110000 ;
			12'h00000973 : data <= 8'b00011000 ;
			12'h00000974 : data <= 8'b00000000 ;
			12'h00000975 : data <= 8'b11001100 ;
			12'h00000976 : data <= 8'b11001100 ;
			12'h00000977 : data <= 8'b11001100 ;
			12'h00000978 : data <= 8'b11001100 ;
			12'h00000979 : data <= 8'b11001100 ;
			12'h0000097A : data <= 8'b11001100 ;
			12'h0000097B : data <= 8'b01110110 ;
			12'h0000097C : data <= 8'b00000000 ;
			12'h0000097D : data <= 8'b00000000 ;
			12'h0000097E : data <= 8'b00000000 ;
			12'h0000097F : data <= 8'b00000000 ;
			12'h00000980 : data <= 8'b00000000 ;
			12'h00000981 : data <= 8'b00000000 ;
			12'h00000982 : data <= 8'b11000110 ;
			12'h00000983 : data <= 8'b00000000 ;
			12'h00000984 : data <= 8'b00000000 ;
			12'h00000985 : data <= 8'b11000110 ;
			12'h00000986 : data <= 8'b11000110 ;
			12'h00000987 : data <= 8'b11000110 ;
			12'h00000988 : data <= 8'b11000110 ;
			12'h00000989 : data <= 8'b11000110 ;
			12'h0000098A : data <= 8'b11000110 ;
			12'h0000098B : data <= 8'b01111110 ;
			12'h0000098C : data <= 8'b00000110 ;
			12'h0000098D : data <= 8'b00001100 ;
			12'h0000098E : data <= 8'b01111000 ;
			12'h0000098F : data <= 8'b00000000 ;
			12'h00000990 : data <= 8'b00000000 ;
			12'h00000991 : data <= 8'b11000110 ;
			12'h00000992 : data <= 8'b00000000 ;
			12'h00000993 : data <= 8'b01111100 ;
			12'h00000994 : data <= 8'b11000110 ;
			12'h00000995 : data <= 8'b11000110 ;
			12'h00000996 : data <= 8'b11000110 ;
			12'h00000997 : data <= 8'b11000110 ;
			12'h00000998 : data <= 8'b11000110 ;
			12'h00000999 : data <= 8'b11000110 ;
			12'h0000099A : data <= 8'b11000110 ;
			12'h0000099B : data <= 8'b01111100 ;
			12'h0000099C : data <= 8'b00000000 ;
			12'h0000099D : data <= 8'b00000000 ;
			12'h0000099E : data <= 8'b00000000 ;
			12'h0000099F : data <= 8'b00000000 ;
			12'h000009A0 : data <= 8'b00000000 ;
			12'h000009A1 : data <= 8'b11000110 ;
			12'h000009A2 : data <= 8'b00000000 ;
			12'h000009A3 : data <= 8'b11000110 ;
			12'h000009A4 : data <= 8'b11000110 ;
			12'h000009A5 : data <= 8'b11000110 ;
			12'h000009A6 : data <= 8'b11000110 ;
			12'h000009A7 : data <= 8'b11000110 ;
			12'h000009A8 : data <= 8'b11000110 ;
			12'h000009A9 : data <= 8'b11000110 ;
			12'h000009AA : data <= 8'b11000110 ;
			12'h000009AB : data <= 8'b01111100 ;
			12'h000009AC : data <= 8'b00000000 ;
			12'h000009AD : data <= 8'b00000000 ;
			12'h000009AE : data <= 8'b00000000 ;
			12'h000009AF : data <= 8'b00000000 ;
			12'h000009B0 : data <= 8'b00000000 ;
			12'h000009B1 : data <= 8'b00011000 ;
			12'h000009B2 : data <= 8'b00011000 ;
			12'h000009B3 : data <= 8'b00111100 ;
			12'h000009B4 : data <= 8'b01100110 ;
			12'h000009B5 : data <= 8'b01100000 ;
			12'h000009B6 : data <= 8'b01100000 ;
			12'h000009B7 : data <= 8'b01100000 ;
			12'h000009B8 : data <= 8'b01100110 ;
			12'h000009B9 : data <= 8'b00111100 ;
			12'h000009BA : data <= 8'b00011000 ;
			12'h000009BB : data <= 8'b00011000 ;
			12'h000009BC : data <= 8'b00000000 ;
			12'h000009BD : data <= 8'b00000000 ;
			12'h000009BE : data <= 8'b00000000 ;
			12'h000009BF : data <= 8'b00000000 ;
			12'h000009C0 : data <= 8'b00000000 ;
			12'h000009C1 : data <= 8'b00111000 ;
			12'h000009C2 : data <= 8'b01101100 ;
			12'h000009C3 : data <= 8'b01100100 ;
			12'h000009C4 : data <= 8'b01100000 ;
			12'h000009C5 : data <= 8'b11110000 ;
			12'h000009C6 : data <= 8'b01100000 ;
			12'h000009C7 : data <= 8'b01100000 ;
			12'h000009C8 : data <= 8'b01100000 ;
			12'h000009C9 : data <= 8'b01100000 ;
			12'h000009CA : data <= 8'b11100110 ;
			12'h000009CB : data <= 8'b11111100 ;
			12'h000009CC : data <= 8'b00000000 ;
			12'h000009CD : data <= 8'b00000000 ;
			12'h000009CE : data <= 8'b00000000 ;
			12'h000009CF : data <= 8'b00000000 ;
			12'h000009D0 : data <= 8'b00000000 ;
			12'h000009D1 : data <= 8'b00000000 ;
			12'h000009D2 : data <= 8'b01100110 ;
			12'h000009D3 : data <= 8'b01100110 ;
			12'h000009D4 : data <= 8'b00111100 ;
			12'h000009D5 : data <= 8'b00011000 ;
			12'h000009D6 : data <= 8'b01111110 ;
			12'h000009D7 : data <= 8'b00011000 ;
			12'h000009D8 : data <= 8'b01111110 ;
			12'h000009D9 : data <= 8'b00011000 ;
			12'h000009DA : data <= 8'b00011000 ;
			12'h000009DB : data <= 8'b00011000 ;
			12'h000009DC : data <= 8'b00000000 ;
			12'h000009DD : data <= 8'b00000000 ;
			12'h000009DE : data <= 8'b00000000 ;
			12'h000009DF : data <= 8'b00000000 ;
			12'h000009E0 : data <= 8'b00000000 ;
			12'h000009E1 : data <= 8'b11111000 ;
			12'h000009E2 : data <= 8'b11001100 ;
			12'h000009E3 : data <= 8'b11001100 ;
			12'h000009E4 : data <= 8'b11111000 ;
			12'h000009E5 : data <= 8'b11000100 ;
			12'h000009E6 : data <= 8'b11001100 ;
			12'h000009E7 : data <= 8'b11011110 ;
			12'h000009E8 : data <= 8'b11001100 ;
			12'h000009E9 : data <= 8'b11001100 ;
			12'h000009EA : data <= 8'b11001100 ;
			12'h000009EB : data <= 8'b11000110 ;
			12'h000009EC : data <= 8'b00000000 ;
			12'h000009ED : data <= 8'b00000000 ;
			12'h000009EE : data <= 8'b00000000 ;
			12'h000009EF : data <= 8'b00000000 ;
			12'h000009F0 : data <= 8'b00000000 ;
			12'h000009F1 : data <= 8'b00001110 ;
			12'h000009F2 : data <= 8'b00011011 ;
			12'h000009F3 : data <= 8'b00011000 ;
			12'h000009F4 : data <= 8'b00011000 ;
			12'h000009F5 : data <= 8'b00011000 ;
			12'h000009F6 : data <= 8'b01111110 ;
			12'h000009F7 : data <= 8'b00011000 ;
			12'h000009F8 : data <= 8'b00011000 ;
			12'h000009F9 : data <= 8'b00011000 ;
			12'h000009FA : data <= 8'b00011000 ;
			12'h000009FB : data <= 8'b00011000 ;
			12'h000009FC : data <= 8'b11011000 ;
			12'h000009FD : data <= 8'b01110000 ;
			12'h000009FE : data <= 8'b00000000 ;
			12'h000009FF : data <= 8'b00000000 ;
			12'h00000A00 : data <= 8'b00000000 ;
			12'h00000A01 : data <= 8'b00011000 ;
			12'h00000A02 : data <= 8'b00110000 ;
			12'h00000A03 : data <= 8'b01100000 ;
			12'h00000A04 : data <= 8'b00000000 ;
			12'h00000A05 : data <= 8'b01111000 ;
			12'h00000A06 : data <= 8'b00001100 ;
			12'h00000A07 : data <= 8'b01111100 ;
			12'h00000A08 : data <= 8'b11001100 ;
			12'h00000A09 : data <= 8'b11001100 ;
			12'h00000A0A : data <= 8'b11001100 ;
			12'h00000A0B : data <= 8'b01110110 ;
			12'h00000A0C : data <= 8'b00000000 ;
			12'h00000A0D : data <= 8'b00000000 ;
			12'h00000A0E : data <= 8'b00000000 ;
			12'h00000A0F : data <= 8'b00000000 ;
			12'h00000A10 : data <= 8'b00000000 ;
			12'h00000A11 : data <= 8'b00001100 ;
			12'h00000A12 : data <= 8'b00011000 ;
			12'h00000A13 : data <= 8'b00110000 ;
			12'h00000A14 : data <= 8'b00000000 ;
			12'h00000A15 : data <= 8'b00111000 ;
			12'h00000A16 : data <= 8'b00011000 ;
			12'h00000A17 : data <= 8'b00011000 ;
			12'h00000A18 : data <= 8'b00011000 ;
			12'h00000A19 : data <= 8'b00011000 ;
			12'h00000A1A : data <= 8'b00011000 ;
			12'h00000A1B : data <= 8'b00111100 ;
			12'h00000A1C : data <= 8'b00000000 ;
			12'h00000A1D : data <= 8'b00000000 ;
			12'h00000A1E : data <= 8'b00000000 ;
			12'h00000A1F : data <= 8'b00000000 ;
			12'h00000A20 : data <= 8'b00000000 ;
			12'h00000A21 : data <= 8'b00011000 ;
			12'h00000A22 : data <= 8'b00110000 ;
			12'h00000A23 : data <= 8'b01100000 ;
			12'h00000A24 : data <= 8'b00000000 ;
			12'h00000A25 : data <= 8'b01111100 ;
			12'h00000A26 : data <= 8'b11000110 ;
			12'h00000A27 : data <= 8'b11000110 ;
			12'h00000A28 : data <= 8'b11000110 ;
			12'h00000A29 : data <= 8'b11000110 ;
			12'h00000A2A : data <= 8'b11000110 ;
			12'h00000A2B : data <= 8'b01111100 ;
			12'h00000A2C : data <= 8'b00000000 ;
			12'h00000A2D : data <= 8'b00000000 ;
			12'h00000A2E : data <= 8'b00000000 ;
			12'h00000A2F : data <= 8'b00000000 ;
			12'h00000A30 : data <= 8'b00000000 ;
			12'h00000A31 : data <= 8'b00011000 ;
			12'h00000A32 : data <= 8'b00110000 ;
			12'h00000A33 : data <= 8'b01100000 ;
			12'h00000A34 : data <= 8'b00000000 ;
			12'h00000A35 : data <= 8'b11001100 ;
			12'h00000A36 : data <= 8'b11001100 ;
			12'h00000A37 : data <= 8'b11001100 ;
			12'h00000A38 : data <= 8'b11001100 ;
			12'h00000A39 : data <= 8'b11001100 ;
			12'h00000A3A : data <= 8'b11001100 ;
			12'h00000A3B : data <= 8'b01110110 ;
			12'h00000A3C : data <= 8'b00000000 ;
			12'h00000A3D : data <= 8'b00000000 ;
			12'h00000A3E : data <= 8'b00000000 ;
			12'h00000A3F : data <= 8'b00000000 ;
			12'h00000A40 : data <= 8'b00000000 ;
			12'h00000A41 : data <= 8'b00000000 ;
			12'h00000A42 : data <= 8'b01110110 ;
			12'h00000A43 : data <= 8'b11011100 ;
			12'h00000A44 : data <= 8'b00000000 ;
			12'h00000A45 : data <= 8'b11011100 ;
			12'h00000A46 : data <= 8'b01100110 ;
			12'h00000A47 : data <= 8'b01100110 ;
			12'h00000A48 : data <= 8'b01100110 ;
			12'h00000A49 : data <= 8'b01100110 ;
			12'h00000A4A : data <= 8'b01100110 ;
			12'h00000A4B : data <= 8'b01100110 ;
			12'h00000A4C : data <= 8'b00000000 ;
			12'h00000A4D : data <= 8'b00000000 ;
			12'h00000A4E : data <= 8'b00000000 ;
			12'h00000A4F : data <= 8'b00000000 ;
			12'h00000A50 : data <= 8'b01110110 ;
			12'h00000A51 : data <= 8'b11011100 ;
			12'h00000A52 : data <= 8'b00000000 ;
			12'h00000A53 : data <= 8'b11000110 ;
			12'h00000A54 : data <= 8'b11100110 ;
			12'h00000A55 : data <= 8'b11110110 ;
			12'h00000A56 : data <= 8'b11111110 ;
			12'h00000A57 : data <= 8'b11011110 ;
			12'h00000A58 : data <= 8'b11001110 ;
			12'h00000A59 : data <= 8'b11000110 ;
			12'h00000A5A : data <= 8'b11000110 ;
			12'h00000A5B : data <= 8'b11000110 ;
			12'h00000A5C : data <= 8'b00000000 ;
			12'h00000A5D : data <= 8'b00000000 ;
			12'h00000A5E : data <= 8'b00000000 ;
			12'h00000A5F : data <= 8'b00000000 ;
			12'h00000A60 : data <= 8'b00000000 ;
			12'h00000A61 : data <= 8'b00111100 ;
			12'h00000A62 : data <= 8'b01101100 ;
			12'h00000A63 : data <= 8'b01101100 ;
			12'h00000A64 : data <= 8'b00111110 ;
			12'h00000A65 : data <= 8'b00000000 ;
			12'h00000A66 : data <= 8'b01111110 ;
			12'h00000A67 : data <= 8'b00000000 ;
			12'h00000A68 : data <= 8'b00000000 ;
			12'h00000A69 : data <= 8'b00000000 ;
			12'h00000A6A : data <= 8'b00000000 ;
			12'h00000A6B : data <= 8'b00000000 ;
			12'h00000A6C : data <= 8'b00000000 ;
			12'h00000A6D : data <= 8'b00000000 ;
			12'h00000A6E : data <= 8'b00000000 ;
			12'h00000A6F : data <= 8'b00000000 ;
			12'h00000A70 : data <= 8'b00000000 ;
			12'h00000A71 : data <= 8'b00111000 ;
			12'h00000A72 : data <= 8'b01101100 ;
			12'h00000A73 : data <= 8'b01101100 ;
			12'h00000A74 : data <= 8'b00111000 ;
			12'h00000A75 : data <= 8'b00000000 ;
			12'h00000A76 : data <= 8'b01111100 ;
			12'h00000A77 : data <= 8'b00000000 ;
			12'h00000A78 : data <= 8'b00000000 ;
			12'h00000A79 : data <= 8'b00000000 ;
			12'h00000A7A : data <= 8'b00000000 ;
			12'h00000A7B : data <= 8'b00000000 ;
			12'h00000A7C : data <= 8'b00000000 ;
			12'h00000A7D : data <= 8'b00000000 ;
			12'h00000A7E : data <= 8'b00000000 ;
			12'h00000A7F : data <= 8'b00000000 ;
			12'h00000A80 : data <= 8'b00000000 ;
			12'h00000A81 : data <= 8'b00000000 ;
			12'h00000A82 : data <= 8'b00110000 ;
			12'h00000A83 : data <= 8'b00110000 ;
			12'h00000A84 : data <= 8'b00000000 ;
			12'h00000A85 : data <= 8'b00110000 ;
			12'h00000A86 : data <= 8'b00110000 ;
			12'h00000A87 : data <= 8'b01100000 ;
			12'h00000A88 : data <= 8'b11000000 ;
			12'h00000A89 : data <= 8'b11000110 ;
			12'h00000A8A : data <= 8'b11000110 ;
			12'h00000A8B : data <= 8'b01111100 ;
			12'h00000A8C : data <= 8'b00000000 ;
			12'h00000A8D : data <= 8'b00000000 ;
			12'h00000A8E : data <= 8'b00000000 ;
			12'h00000A8F : data <= 8'b00000000 ;
			12'h00000A90 : data <= 8'b00000000 ;
			12'h00000A91 : data <= 8'b00000000 ;
			12'h00000A92 : data <= 8'b00000000 ;
			12'h00000A93 : data <= 8'b00000000 ;
			12'h00000A94 : data <= 8'b00000000 ;
			12'h00000A95 : data <= 8'b00000000 ;
			12'h00000A96 : data <= 8'b11111110 ;
			12'h00000A97 : data <= 8'b11000000 ;
			12'h00000A98 : data <= 8'b11000000 ;
			12'h00000A99 : data <= 8'b11000000 ;
			12'h00000A9A : data <= 8'b11000000 ;
			12'h00000A9B : data <= 8'b00000000 ;
			12'h00000A9C : data <= 8'b00000000 ;
			12'h00000A9D : data <= 8'b00000000 ;
			12'h00000A9E : data <= 8'b00000000 ;
			12'h00000A9F : data <= 8'b00000000 ;
			12'h00000AA0 : data <= 8'b00000000 ;
			12'h00000AA1 : data <= 8'b00000000 ;
			12'h00000AA2 : data <= 8'b00000000 ;
			12'h00000AA3 : data <= 8'b00000000 ;
			12'h00000AA4 : data <= 8'b00000000 ;
			12'h00000AA5 : data <= 8'b00000000 ;
			12'h00000AA6 : data <= 8'b11111110 ;
			12'h00000AA7 : data <= 8'b00000110 ;
			12'h00000AA8 : data <= 8'b00000110 ;
			12'h00000AA9 : data <= 8'b00000110 ;
			12'h00000AAA : data <= 8'b00000110 ;
			12'h00000AAB : data <= 8'b00000000 ;
			12'h00000AAC : data <= 8'b00000000 ;
			12'h00000AAD : data <= 8'b00000000 ;
			12'h00000AAE : data <= 8'b00000000 ;
			12'h00000AAF : data <= 8'b00000000 ;
			12'h00000AB0 : data <= 8'b00000000 ;
			12'h00000AB1 : data <= 8'b11000000 ;
			12'h00000AB2 : data <= 8'b11000000 ;
			12'h00000AB3 : data <= 8'b11000010 ;
			12'h00000AB4 : data <= 8'b11000110 ;
			12'h00000AB5 : data <= 8'b11001100 ;
			12'h00000AB6 : data <= 8'b00011000 ;
			12'h00000AB7 : data <= 8'b00110000 ;
			12'h00000AB8 : data <= 8'b01100000 ;
			12'h00000AB9 : data <= 8'b11011100 ;
			12'h00000ABA : data <= 8'b10000110 ;
			12'h00000ABB : data <= 8'b00001100 ;
			12'h00000ABC : data <= 8'b00011000 ;
			12'h00000ABD : data <= 8'b00111110 ;
			12'h00000ABE : data <= 8'b00000000 ;
			12'h00000ABF : data <= 8'b00000000 ;
			12'h00000AC0 : data <= 8'b00000000 ;
			12'h00000AC1 : data <= 8'b11000000 ;
			12'h00000AC2 : data <= 8'b11000000 ;
			12'h00000AC3 : data <= 8'b11000010 ;
			12'h00000AC4 : data <= 8'b11000110 ;
			12'h00000AC5 : data <= 8'b11001100 ;
			12'h00000AC6 : data <= 8'b00011000 ;
			12'h00000AC7 : data <= 8'b00110000 ;
			12'h00000AC8 : data <= 8'b01100110 ;
			12'h00000AC9 : data <= 8'b11001110 ;
			12'h00000ACA : data <= 8'b10011110 ;
			12'h00000ACB : data <= 8'b00111110 ;
			12'h00000ACC : data <= 8'b00000110 ;
			12'h00000ACD : data <= 8'b00000110 ;
			12'h00000ACE : data <= 8'b00000000 ;
			12'h00000ACF : data <= 8'b00000000 ;
			12'h00000AD0 : data <= 8'b00000000 ;
			12'h00000AD1 : data <= 8'b00000000 ;
			12'h00000AD2 : data <= 8'b00011000 ;
			12'h00000AD3 : data <= 8'b00011000 ;
			12'h00000AD4 : data <= 8'b00000000 ;
			12'h00000AD5 : data <= 8'b00011000 ;
			12'h00000AD6 : data <= 8'b00011000 ;
			12'h00000AD7 : data <= 8'b00011000 ;
			12'h00000AD8 : data <= 8'b00111100 ;
			12'h00000AD9 : data <= 8'b00111100 ;
			12'h00000ADA : data <= 8'b00111100 ;
			12'h00000ADB : data <= 8'b00011000 ;
			12'h00000ADC : data <= 8'b00000000 ;
			12'h00000ADD : data <= 8'b00000000 ;
			12'h00000ADE : data <= 8'b00000000 ;
			12'h00000ADF : data <= 8'b00000000 ;
			12'h00000AE0 : data <= 8'b00000000 ;
			12'h00000AE1 : data <= 8'b00000000 ;
			12'h00000AE2 : data <= 8'b00000000 ;
			12'h00000AE3 : data <= 8'b00000000 ;
			12'h00000AE4 : data <= 8'b00000000 ;
			12'h00000AE5 : data <= 8'b00110110 ;
			12'h00000AE6 : data <= 8'b01101100 ;
			12'h00000AE7 : data <= 8'b11011000 ;
			12'h00000AE8 : data <= 8'b01101100 ;
			12'h00000AE9 : data <= 8'b00110110 ;
			12'h00000AEA : data <= 8'b00000000 ;
			12'h00000AEB : data <= 8'b00000000 ;
			12'h00000AEC : data <= 8'b00000000 ;
			12'h00000AED : data <= 8'b00000000 ;
			12'h00000AEE : data <= 8'b00000000 ;
			12'h00000AEF : data <= 8'b00000000 ;
			12'h00000AF0 : data <= 8'b00000000 ;
			12'h00000AF1 : data <= 8'b00000000 ;
			12'h00000AF2 : data <= 8'b00000000 ;
			12'h00000AF3 : data <= 8'b00000000 ;
			12'h00000AF4 : data <= 8'b00000000 ;
			12'h00000AF5 : data <= 8'b11011000 ;
			12'h00000AF6 : data <= 8'b01101100 ;
			12'h00000AF7 : data <= 8'b00110110 ;
			12'h00000AF8 : data <= 8'b01101100 ;
			12'h00000AF9 : data <= 8'b11011000 ;
			12'h00000AFA : data <= 8'b00000000 ;
			12'h00000AFB : data <= 8'b00000000 ;
			12'h00000AFC : data <= 8'b00000000 ;
			12'h00000AFD : data <= 8'b00000000 ;
			12'h00000AFE : data <= 8'b00000000 ;
			12'h00000AFF : data <= 8'b00000000 ;
			12'h00000B00 : data <= 8'b00010001 ;
			12'h00000B01 : data <= 8'b01000100 ;
			12'h00000B02 : data <= 8'b00010001 ;
			12'h00000B03 : data <= 8'b01000100 ;
			12'h00000B04 : data <= 8'b00010001 ;
			12'h00000B05 : data <= 8'b01000100 ;
			12'h00000B06 : data <= 8'b00010001 ;
			12'h00000B07 : data <= 8'b01000100 ;
			12'h00000B08 : data <= 8'b00010001 ;
			12'h00000B09 : data <= 8'b01000100 ;
			12'h00000B0A : data <= 8'b00010001 ;
			12'h00000B0B : data <= 8'b01000100 ;
			12'h00000B0C : data <= 8'b00010001 ;
			12'h00000B0D : data <= 8'b01000100 ;
			12'h00000B0E : data <= 8'b00010001 ;
			12'h00000B0F : data <= 8'b01000100 ;
			12'h00000B10 : data <= 8'b01010101 ;
			12'h00000B11 : data <= 8'b10101010 ;
			12'h00000B12 : data <= 8'b01010101 ;
			12'h00000B13 : data <= 8'b10101010 ;
			12'h00000B14 : data <= 8'b01010101 ;
			12'h00000B15 : data <= 8'b10101010 ;
			12'h00000B16 : data <= 8'b01010101 ;
			12'h00000B17 : data <= 8'b10101010 ;
			12'h00000B18 : data <= 8'b01010101 ;
			12'h00000B19 : data <= 8'b10101010 ;
			12'h00000B1A : data <= 8'b01010101 ;
			12'h00000B1B : data <= 8'b10101010 ;
			12'h00000B1C : data <= 8'b01010101 ;
			12'h00000B1D : data <= 8'b10101010 ;
			12'h00000B1E : data <= 8'b01010101 ;
			12'h00000B1F : data <= 8'b10101010 ;
			12'h00000B20 : data <= 8'b11011101 ;
			12'h00000B21 : data <= 8'b01110111 ;
			12'h00000B22 : data <= 8'b11011101 ;
			12'h00000B23 : data <= 8'b01110111 ;
			12'h00000B24 : data <= 8'b11011101 ;
			12'h00000B25 : data <= 8'b01110111 ;
			12'h00000B26 : data <= 8'b11011101 ;
			12'h00000B27 : data <= 8'b01110111 ;
			12'h00000B28 : data <= 8'b11011101 ;
			12'h00000B29 : data <= 8'b01110111 ;
			12'h00000B2A : data <= 8'b11011101 ;
			12'h00000B2B : data <= 8'b01110111 ;
			12'h00000B2C : data <= 8'b11011101 ;
			12'h00000B2D : data <= 8'b01110111 ;
			12'h00000B2E : data <= 8'b11011101 ;
			12'h00000B2F : data <= 8'b01110111 ;
			12'h00000B30 : data <= 8'b00011000 ;
			12'h00000B31 : data <= 8'b00011000 ;
			12'h00000B32 : data <= 8'b00011000 ;
			12'h00000B33 : data <= 8'b00011000 ;
			12'h00000B34 : data <= 8'b00011000 ;
			12'h00000B35 : data <= 8'b00011000 ;
			12'h00000B36 : data <= 8'b00011000 ;
			12'h00000B37 : data <= 8'b00011000 ;
			12'h00000B38 : data <= 8'b00011000 ;
			12'h00000B39 : data <= 8'b00011000 ;
			12'h00000B3A : data <= 8'b00011000 ;
			12'h00000B3B : data <= 8'b00011000 ;
			12'h00000B3C : data <= 8'b00011000 ;
			12'h00000B3D : data <= 8'b00011000 ;
			12'h00000B3E : data <= 8'b00011000 ;
			12'h00000B3F : data <= 8'b00011000 ;
			12'h00000B40 : data <= 8'b00011000 ;
			12'h00000B41 : data <= 8'b00011000 ;
			12'h00000B42 : data <= 8'b00011000 ;
			12'h00000B43 : data <= 8'b00011000 ;
			12'h00000B44 : data <= 8'b00011000 ;
			12'h00000B45 : data <= 8'b00011000 ;
			12'h00000B46 : data <= 8'b00011000 ;
			12'h00000B47 : data <= 8'b11111000 ;
			12'h00000B48 : data <= 8'b00011000 ;
			12'h00000B49 : data <= 8'b00011000 ;
			12'h00000B4A : data <= 8'b00011000 ;
			12'h00000B4B : data <= 8'b00011000 ;
			12'h00000B4C : data <= 8'b00011000 ;
			12'h00000B4D : data <= 8'b00011000 ;
			12'h00000B4E : data <= 8'b00011000 ;
			12'h00000B4F : data <= 8'b00011000 ;
			12'h00000B50 : data <= 8'b00011000 ;
			12'h00000B51 : data <= 8'b00011000 ;
			12'h00000B52 : data <= 8'b00011000 ;
			12'h00000B53 : data <= 8'b00011000 ;
			12'h00000B54 : data <= 8'b00011000 ;
			12'h00000B55 : data <= 8'b11111000 ;
			12'h00000B56 : data <= 8'b00011000 ;
			12'h00000B57 : data <= 8'b11111000 ;
			12'h00000B58 : data <= 8'b00011000 ;
			12'h00000B59 : data <= 8'b00011000 ;
			12'h00000B5A : data <= 8'b00011000 ;
			12'h00000B5B : data <= 8'b00011000 ;
			12'h00000B5C : data <= 8'b00011000 ;
			12'h00000B5D : data <= 8'b00011000 ;
			12'h00000B5E : data <= 8'b00011000 ;
			12'h00000B5F : data <= 8'b00011000 ;
			12'h00000B60 : data <= 8'b00110110 ;
			12'h00000B61 : data <= 8'b00110110 ;
			12'h00000B62 : data <= 8'b00110110 ;
			12'h00000B63 : data <= 8'b00110110 ;
			12'h00000B64 : data <= 8'b00110110 ;
			12'h00000B65 : data <= 8'b00110110 ;
			12'h00000B66 : data <= 8'b00110110 ;
			12'h00000B67 : data <= 8'b11110110 ;
			12'h00000B68 : data <= 8'b00110110 ;
			12'h00000B69 : data <= 8'b00110110 ;
			12'h00000B6A : data <= 8'b00110110 ;
			12'h00000B6B : data <= 8'b00110110 ;
			12'h00000B6C : data <= 8'b00110110 ;
			12'h00000B6D : data <= 8'b00110110 ;
			12'h00000B6E : data <= 8'b00110110 ;
			12'h00000B6F : data <= 8'b00110110 ;
			12'h00000B70 : data <= 8'b00000000 ;
			12'h00000B71 : data <= 8'b00000000 ;
			12'h00000B72 : data <= 8'b00000000 ;
			12'h00000B73 : data <= 8'b00000000 ;
			12'h00000B74 : data <= 8'b00000000 ;
			12'h00000B75 : data <= 8'b00000000 ;
			12'h00000B76 : data <= 8'b00000000 ;
			12'h00000B77 : data <= 8'b11111110 ;
			12'h00000B78 : data <= 8'b00110110 ;
			12'h00000B79 : data <= 8'b00110110 ;
			12'h00000B7A : data <= 8'b00110110 ;
			12'h00000B7B : data <= 8'b00110110 ;
			12'h00000B7C : data <= 8'b00110110 ;
			12'h00000B7D : data <= 8'b00110110 ;
			12'h00000B7E : data <= 8'b00110110 ;
			12'h00000B7F : data <= 8'b00110110 ;
			12'h00000B80 : data <= 8'b00000000 ;
			12'h00000B81 : data <= 8'b00000000 ;
			12'h00000B82 : data <= 8'b00000000 ;
			12'h00000B83 : data <= 8'b00000000 ;
			12'h00000B84 : data <= 8'b00000000 ;
			12'h00000B85 : data <= 8'b11111000 ;
			12'h00000B86 : data <= 8'b00011000 ;
			12'h00000B87 : data <= 8'b11111000 ;
			12'h00000B88 : data <= 8'b00011000 ;
			12'h00000B89 : data <= 8'b00011000 ;
			12'h00000B8A : data <= 8'b00011000 ;
			12'h00000B8B : data <= 8'b00011000 ;
			12'h00000B8C : data <= 8'b00011000 ;
			12'h00000B8D : data <= 8'b00011000 ;
			12'h00000B8E : data <= 8'b00011000 ;
			12'h00000B8F : data <= 8'b00011000 ;
			12'h00000B90 : data <= 8'b00110110 ;
			12'h00000B91 : data <= 8'b00110110 ;
			12'h00000B92 : data <= 8'b00110110 ;
			12'h00000B93 : data <= 8'b00110110 ;
			12'h00000B94 : data <= 8'b00110110 ;
			12'h00000B95 : data <= 8'b11110110 ;
			12'h00000B96 : data <= 8'b00000110 ;
			12'h00000B97 : data <= 8'b11110110 ;
			12'h00000B98 : data <= 8'b00110110 ;
			12'h00000B99 : data <= 8'b00110110 ;
			12'h00000B9A : data <= 8'b00110110 ;
			12'h00000B9B : data <= 8'b00110110 ;
			12'h00000B9C : data <= 8'b00110110 ;
			12'h00000B9D : data <= 8'b00110110 ;
			12'h00000B9E : data <= 8'b00110110 ;
			12'h00000B9F : data <= 8'b00110110 ;
			12'h00000BA0 : data <= 8'b00110110 ;
			12'h00000BA1 : data <= 8'b00110110 ;
			12'h00000BA2 : data <= 8'b00110110 ;
			12'h00000BA3 : data <= 8'b00110110 ;
			12'h00000BA4 : data <= 8'b00110110 ;
			12'h00000BA5 : data <= 8'b00110110 ;
			12'h00000BA6 : data <= 8'b00110110 ;
			12'h00000BA7 : data <= 8'b00110110 ;
			12'h00000BA8 : data <= 8'b00110110 ;
			12'h00000BA9 : data <= 8'b00110110 ;
			12'h00000BAA : data <= 8'b00110110 ;
			12'h00000BAB : data <= 8'b00110110 ;
			12'h00000BAC : data <= 8'b00110110 ;
			12'h00000BAD : data <= 8'b00110110 ;
			12'h00000BAE : data <= 8'b00110110 ;
			12'h00000BAF : data <= 8'b00110110 ;
			12'h00000BB0 : data <= 8'b00000000 ;
			12'h00000BB1 : data <= 8'b00000000 ;
			12'h00000BB2 : data <= 8'b00000000 ;
			12'h00000BB3 : data <= 8'b00000000 ;
			12'h00000BB4 : data <= 8'b00000000 ;
			12'h00000BB5 : data <= 8'b11111110 ;
			12'h00000BB6 : data <= 8'b00000110 ;
			12'h00000BB7 : data <= 8'b11110110 ;
			12'h00000BB8 : data <= 8'b00110110 ;
			12'h00000BB9 : data <= 8'b00110110 ;
			12'h00000BBA : data <= 8'b00110110 ;
			12'h00000BBB : data <= 8'b00110110 ;
			12'h00000BBC : data <= 8'b00110110 ;
			12'h00000BBD : data <= 8'b00110110 ;
			12'h00000BBE : data <= 8'b00110110 ;
			12'h00000BBF : data <= 8'b00110110 ;
			12'h00000BC0 : data <= 8'b00110110 ;
			12'h00000BC1 : data <= 8'b00110110 ;
			12'h00000BC2 : data <= 8'b00110110 ;
			12'h00000BC3 : data <= 8'b00110110 ;
			12'h00000BC4 : data <= 8'b00110110 ;
			12'h00000BC5 : data <= 8'b11110110 ;
			12'h00000BC6 : data <= 8'b00000110 ;
			12'h00000BC7 : data <= 8'b11111110 ;
			12'h00000BC8 : data <= 8'b00000000 ;
			12'h00000BC9 : data <= 8'b00000000 ;
			12'h00000BCA : data <= 8'b00000000 ;
			12'h00000BCB : data <= 8'b00000000 ;
			12'h00000BCC : data <= 8'b00000000 ;
			12'h00000BCD : data <= 8'b00000000 ;
			12'h00000BCE : data <= 8'b00000000 ;
			12'h00000BCF : data <= 8'b00000000 ;
			12'h00000BD0 : data <= 8'b00110110 ;
			12'h00000BD1 : data <= 8'b00110110 ;
			12'h00000BD2 : data <= 8'b00110110 ;
			12'h00000BD3 : data <= 8'b00110110 ;
			12'h00000BD4 : data <= 8'b00110110 ;
			12'h00000BD5 : data <= 8'b00110110 ;
			12'h00000BD6 : data <= 8'b00110110 ;
			12'h00000BD7 : data <= 8'b11111110 ;
			12'h00000BD8 : data <= 8'b00000000 ;
			12'h00000BD9 : data <= 8'b00000000 ;
			12'h00000BDA : data <= 8'b00000000 ;
			12'h00000BDB : data <= 8'b00000000 ;
			12'h00000BDC : data <= 8'b00000000 ;
			12'h00000BDD : data <= 8'b00000000 ;
			12'h00000BDE : data <= 8'b00000000 ;
			12'h00000BDF : data <= 8'b00000000 ;
			12'h00000BE0 : data <= 8'b00011000 ;
			12'h00000BE1 : data <= 8'b00011000 ;
			12'h00000BE2 : data <= 8'b00011000 ;
			12'h00000BE3 : data <= 8'b00011000 ;
			12'h00000BE4 : data <= 8'b00011000 ;
			12'h00000BE5 : data <= 8'b11111000 ;
			12'h00000BE6 : data <= 8'b00011000 ;
			12'h00000BE7 : data <= 8'b11111000 ;
			12'h00000BE8 : data <= 8'b00000000 ;
			12'h00000BE9 : data <= 8'b00000000 ;
			12'h00000BEA : data <= 8'b00000000 ;
			12'h00000BEB : data <= 8'b00000000 ;
			12'h00000BEC : data <= 8'b00000000 ;
			12'h00000BED : data <= 8'b00000000 ;
			12'h00000BEE : data <= 8'b00000000 ;
			12'h00000BEF : data <= 8'b00000000 ;
			12'h00000BF0 : data <= 8'b00000000 ;
			12'h00000BF1 : data <= 8'b00000000 ;
			12'h00000BF2 : data <= 8'b00000000 ;
			12'h00000BF3 : data <= 8'b00000000 ;
			12'h00000BF4 : data <= 8'b00000000 ;
			12'h00000BF5 : data <= 8'b00000000 ;
			12'h00000BF6 : data <= 8'b00000000 ;
			12'h00000BF7 : data <= 8'b11111000 ;
			12'h00000BF8 : data <= 8'b00011000 ;
			12'h00000BF9 : data <= 8'b00011000 ;
			12'h00000BFA : data <= 8'b00011000 ;
			12'h00000BFB : data <= 8'b00011000 ;
			12'h00000BFC : data <= 8'b00011000 ;
			12'h00000BFD : data <= 8'b00011000 ;
			12'h00000BFE : data <= 8'b00011000 ;
			12'h00000BFF : data <= 8'b00011000 ;
			12'h00000C00 : data <= 8'b00011000 ;
			12'h00000C01 : data <= 8'b00011000 ;
			12'h00000C02 : data <= 8'b00011000 ;
			12'h00000C03 : data <= 8'b00011000 ;
			12'h00000C04 : data <= 8'b00011000 ;
			12'h00000C05 : data <= 8'b00011000 ;
			12'h00000C06 : data <= 8'b00011000 ;
			12'h00000C07 : data <= 8'b00011111 ;
			12'h00000C08 : data <= 8'b00000000 ;
			12'h00000C09 : data <= 8'b00000000 ;
			12'h00000C0A : data <= 8'b00000000 ;
			12'h00000C0B : data <= 8'b00000000 ;
			12'h00000C0C : data <= 8'b00000000 ;
			12'h00000C0D : data <= 8'b00000000 ;
			12'h00000C0E : data <= 8'b00000000 ;
			12'h00000C0F : data <= 8'b00000000 ;
			12'h00000C10 : data <= 8'b00011000 ;
			12'h00000C11 : data <= 8'b00011000 ;
			12'h00000C12 : data <= 8'b00011000 ;
			12'h00000C13 : data <= 8'b00011000 ;
			12'h00000C14 : data <= 8'b00011000 ;
			12'h00000C15 : data <= 8'b00011000 ;
			12'h00000C16 : data <= 8'b00011000 ;
			12'h00000C17 : data <= 8'b11111111 ;
			12'h00000C18 : data <= 8'b00000000 ;
			12'h00000C19 : data <= 8'b00000000 ;
			12'h00000C1A : data <= 8'b00000000 ;
			12'h00000C1B : data <= 8'b00000000 ;
			12'h00000C1C : data <= 8'b00000000 ;
			12'h00000C1D : data <= 8'b00000000 ;
			12'h00000C1E : data <= 8'b00000000 ;
			12'h00000C1F : data <= 8'b00000000 ;
			12'h00000C20 : data <= 8'b00000000 ;
			12'h00000C21 : data <= 8'b00000000 ;
			12'h00000C22 : data <= 8'b00000000 ;
			12'h00000C23 : data <= 8'b00000000 ;
			12'h00000C24 : data <= 8'b00000000 ;
			12'h00000C25 : data <= 8'b00000000 ;
			12'h00000C26 : data <= 8'b00000000 ;
			12'h00000C27 : data <= 8'b11111111 ;
			12'h00000C28 : data <= 8'b00011000 ;
			12'h00000C29 : data <= 8'b00011000 ;
			12'h00000C2A : data <= 8'b00011000 ;
			12'h00000C2B : data <= 8'b00011000 ;
			12'h00000C2C : data <= 8'b00011000 ;
			12'h00000C2D : data <= 8'b00011000 ;
			12'h00000C2E : data <= 8'b00011000 ;
			12'h00000C2F : data <= 8'b00011000 ;
			12'h00000C30 : data <= 8'b00011000 ;
			12'h00000C31 : data <= 8'b00011000 ;
			12'h00000C32 : data <= 8'b00011000 ;
			12'h00000C33 : data <= 8'b00011000 ;
			12'h00000C34 : data <= 8'b00011000 ;
			12'h00000C35 : data <= 8'b00011000 ;
			12'h00000C36 : data <= 8'b00011000 ;
			12'h00000C37 : data <= 8'b00011111 ;
			12'h00000C38 : data <= 8'b00011000 ;
			12'h00000C39 : data <= 8'b00011000 ;
			12'h00000C3A : data <= 8'b00011000 ;
			12'h00000C3B : data <= 8'b00011000 ;
			12'h00000C3C : data <= 8'b00011000 ;
			12'h00000C3D : data <= 8'b00011000 ;
			12'h00000C3E : data <= 8'b00011000 ;
			12'h00000C3F : data <= 8'b00011000 ;
			12'h00000C40 : data <= 8'b00000000 ;
			12'h00000C41 : data <= 8'b00000000 ;
			12'h00000C42 : data <= 8'b00000000 ;
			12'h00000C43 : data <= 8'b00000000 ;
			12'h00000C44 : data <= 8'b00000000 ;
			12'h00000C45 : data <= 8'b00000000 ;
			12'h00000C46 : data <= 8'b00000000 ;
			12'h00000C47 : data <= 8'b11111111 ;
			12'h00000C48 : data <= 8'b00000000 ;
			12'h00000C49 : data <= 8'b00000000 ;
			12'h00000C4A : data <= 8'b00000000 ;
			12'h00000C4B : data <= 8'b00000000 ;
			12'h00000C4C : data <= 8'b00000000 ;
			12'h00000C4D : data <= 8'b00000000 ;
			12'h00000C4E : data <= 8'b00000000 ;
			12'h00000C4F : data <= 8'b00000000 ;
			12'h00000C50 : data <= 8'b00011000 ;
			12'h00000C51 : data <= 8'b00011000 ;
			12'h00000C52 : data <= 8'b00011000 ;
			12'h00000C53 : data <= 8'b00011000 ;
			12'h00000C54 : data <= 8'b00011000 ;
			12'h00000C55 : data <= 8'b00011000 ;
			12'h00000C56 : data <= 8'b00011000 ;
			12'h00000C57 : data <= 8'b11111111 ;
			12'h00000C58 : data <= 8'b00011000 ;
			12'h00000C59 : data <= 8'b00011000 ;
			12'h00000C5A : data <= 8'b00011000 ;
			12'h00000C5B : data <= 8'b00011000 ;
			12'h00000C5C : data <= 8'b00011000 ;
			12'h00000C5D : data <= 8'b00011000 ;
			12'h00000C5E : data <= 8'b00011000 ;
			12'h00000C5F : data <= 8'b00011000 ;
			12'h00000C60 : data <= 8'b00011000 ;
			12'h00000C61 : data <= 8'b00011000 ;
			12'h00000C62 : data <= 8'b00011000 ;
			12'h00000C63 : data <= 8'b00011000 ;
			12'h00000C64 : data <= 8'b00011000 ;
			12'h00000C65 : data <= 8'b00011111 ;
			12'h00000C66 : data <= 8'b00011000 ;
			12'h00000C67 : data <= 8'b00011111 ;
			12'h00000C68 : data <= 8'b00011000 ;
			12'h00000C69 : data <= 8'b00011000 ;
			12'h00000C6A : data <= 8'b00011000 ;
			12'h00000C6B : data <= 8'b00011000 ;
			12'h00000C6C : data <= 8'b00011000 ;
			12'h00000C6D : data <= 8'b00011000 ;
			12'h00000C6E : data <= 8'b00011000 ;
			12'h00000C6F : data <= 8'b00011000 ;
			12'h00000C70 : data <= 8'b00110110 ;
			12'h00000C71 : data <= 8'b00110110 ;
			12'h00000C72 : data <= 8'b00110110 ;
			12'h00000C73 : data <= 8'b00110110 ;
			12'h00000C74 : data <= 8'b00110110 ;
			12'h00000C75 : data <= 8'b00110110 ;
			12'h00000C76 : data <= 8'b00110110 ;
			12'h00000C77 : data <= 8'b00110111 ;
			12'h00000C78 : data <= 8'b00110110 ;
			12'h00000C79 : data <= 8'b00110110 ;
			12'h00000C7A : data <= 8'b00110110 ;
			12'h00000C7B : data <= 8'b00110110 ;
			12'h00000C7C : data <= 8'b00110110 ;
			12'h00000C7D : data <= 8'b00110110 ;
			12'h00000C7E : data <= 8'b00110110 ;
			12'h00000C7F : data <= 8'b00110110 ;
			12'h00000C80 : data <= 8'b00110110 ;
			12'h00000C81 : data <= 8'b00110110 ;
			12'h00000C82 : data <= 8'b00110110 ;
			12'h00000C83 : data <= 8'b00110110 ;
			12'h00000C84 : data <= 8'b00110110 ;
			12'h00000C85 : data <= 8'b00110111 ;
			12'h00000C86 : data <= 8'b00110000 ;
			12'h00000C87 : data <= 8'b00111111 ;
			12'h00000C88 : data <= 8'b00000000 ;
			12'h00000C89 : data <= 8'b00000000 ;
			12'h00000C8A : data <= 8'b00000000 ;
			12'h00000C8B : data <= 8'b00000000 ;
			12'h00000C8C : data <= 8'b00000000 ;
			12'h00000C8D : data <= 8'b00000000 ;
			12'h00000C8E : data <= 8'b00000000 ;
			12'h00000C8F : data <= 8'b00000000 ;
			12'h00000C90 : data <= 8'b00000000 ;
			12'h00000C91 : data <= 8'b00000000 ;
			12'h00000C92 : data <= 8'b00000000 ;
			12'h00000C93 : data <= 8'b00000000 ;
			12'h00000C94 : data <= 8'b00000000 ;
			12'h00000C95 : data <= 8'b00111111 ;
			12'h00000C96 : data <= 8'b00110000 ;
			12'h00000C97 : data <= 8'b00110111 ;
			12'h00000C98 : data <= 8'b00110110 ;
			12'h00000C99 : data <= 8'b00110110 ;
			12'h00000C9A : data <= 8'b00110110 ;
			12'h00000C9B : data <= 8'b00110110 ;
			12'h00000C9C : data <= 8'b00110110 ;
			12'h00000C9D : data <= 8'b00110110 ;
			12'h00000C9E : data <= 8'b00110110 ;
			12'h00000C9F : data <= 8'b00110110 ;
			12'h00000CA0 : data <= 8'b00110110 ;
			12'h00000CA1 : data <= 8'b00110110 ;
			12'h00000CA2 : data <= 8'b00110110 ;
			12'h00000CA3 : data <= 8'b00110110 ;
			12'h00000CA4 : data <= 8'b00110110 ;
			12'h00000CA5 : data <= 8'b11110111 ;
			12'h00000CA6 : data <= 8'b00000000 ;
			12'h00000CA7 : data <= 8'b11111111 ;
			12'h00000CA8 : data <= 8'b00000000 ;
			12'h00000CA9 : data <= 8'b00000000 ;
			12'h00000CAA : data <= 8'b00000000 ;
			12'h00000CAB : data <= 8'b00000000 ;
			12'h00000CAC : data <= 8'b00000000 ;
			12'h00000CAD : data <= 8'b00000000 ;
			12'h00000CAE : data <= 8'b00000000 ;
			12'h00000CAF : data <= 8'b00000000 ;
			12'h00000CB0 : data <= 8'b00000000 ;
			12'h00000CB1 : data <= 8'b00000000 ;
			12'h00000CB2 : data <= 8'b00000000 ;
			12'h00000CB3 : data <= 8'b00000000 ;
			12'h00000CB4 : data <= 8'b00000000 ;
			12'h00000CB5 : data <= 8'b11111111 ;
			12'h00000CB6 : data <= 8'b00000000 ;
			12'h00000CB7 : data <= 8'b11110111 ;
			12'h00000CB8 : data <= 8'b00110110 ;
			12'h00000CB9 : data <= 8'b00110110 ;
			12'h00000CBA : data <= 8'b00110110 ;
			12'h00000CBB : data <= 8'b00110110 ;
			12'h00000CBC : data <= 8'b00110110 ;
			12'h00000CBD : data <= 8'b00110110 ;
			12'h00000CBE : data <= 8'b00110110 ;
			12'h00000CBF : data <= 8'b00110110 ;
			12'h00000CC0 : data <= 8'b00110110 ;
			12'h00000CC1 : data <= 8'b00110110 ;
			12'h00000CC2 : data <= 8'b00110110 ;
			12'h00000CC3 : data <= 8'b00110110 ;
			12'h00000CC4 : data <= 8'b00110110 ;
			12'h00000CC5 : data <= 8'b00110111 ;
			12'h00000CC6 : data <= 8'b00110000 ;
			12'h00000CC7 : data <= 8'b00110111 ;
			12'h00000CC8 : data <= 8'b00110110 ;
			12'h00000CC9 : data <= 8'b00110110 ;
			12'h00000CCA : data <= 8'b00110110 ;
			12'h00000CCB : data <= 8'b00110110 ;
			12'h00000CCC : data <= 8'b00110110 ;
			12'h00000CCD : data <= 8'b00110110 ;
			12'h00000CCE : data <= 8'b00110110 ;
			12'h00000CCF : data <= 8'b00110110 ;
			12'h00000CD0 : data <= 8'b00000000 ;
			12'h00000CD1 : data <= 8'b00000000 ;
			12'h00000CD2 : data <= 8'b00000000 ;
			12'h00000CD3 : data <= 8'b00000000 ;
			12'h00000CD4 : data <= 8'b00000000 ;
			12'h00000CD5 : data <= 8'b11111111 ;
			12'h00000CD6 : data <= 8'b00000000 ;
			12'h00000CD7 : data <= 8'b11111111 ;
			12'h00000CD8 : data <= 8'b00000000 ;
			12'h00000CD9 : data <= 8'b00000000 ;
			12'h00000CDA : data <= 8'b00000000 ;
			12'h00000CDB : data <= 8'b00000000 ;
			12'h00000CDC : data <= 8'b00000000 ;
			12'h00000CDD : data <= 8'b00000000 ;
			12'h00000CDE : data <= 8'b00000000 ;
			12'h00000CDF : data <= 8'b00000000 ;
			12'h00000CE0 : data <= 8'b00110110 ;
			12'h00000CE1 : data <= 8'b00110110 ;
			12'h00000CE2 : data <= 8'b00110110 ;
			12'h00000CE3 : data <= 8'b00110110 ;
			12'h00000CE4 : data <= 8'b00110110 ;
			12'h00000CE5 : data <= 8'b11110111 ;
			12'h00000CE6 : data <= 8'b00000000 ;
			12'h00000CE7 : data <= 8'b11110111 ;
			12'h00000CE8 : data <= 8'b00110110 ;
			12'h00000CE9 : data <= 8'b00110110 ;
			12'h00000CEA : data <= 8'b00110110 ;
			12'h00000CEB : data <= 8'b00110110 ;
			12'h00000CEC : data <= 8'b00110110 ;
			12'h00000CED : data <= 8'b00110110 ;
			12'h00000CEE : data <= 8'b00110110 ;
			12'h00000CEF : data <= 8'b00110110 ;
			12'h00000CF0 : data <= 8'b00011000 ;
			12'h00000CF1 : data <= 8'b00011000 ;
			12'h00000CF2 : data <= 8'b00011000 ;
			12'h00000CF3 : data <= 8'b00011000 ;
			12'h00000CF4 : data <= 8'b00011000 ;
			12'h00000CF5 : data <= 8'b11111111 ;
			12'h00000CF6 : data <= 8'b00000000 ;
			12'h00000CF7 : data <= 8'b11111111 ;
			12'h00000CF8 : data <= 8'b00000000 ;
			12'h00000CF9 : data <= 8'b00000000 ;
			12'h00000CFA : data <= 8'b00000000 ;
			12'h00000CFB : data <= 8'b00000000 ;
			12'h00000CFC : data <= 8'b00000000 ;
			12'h00000CFD : data <= 8'b00000000 ;
			12'h00000CFE : data <= 8'b00000000 ;
			12'h00000CFF : data <= 8'b00000000 ;
			12'h00000D00 : data <= 8'b00110110 ;
			12'h00000D01 : data <= 8'b00110110 ;
			12'h00000D02 : data <= 8'b00110110 ;
			12'h00000D03 : data <= 8'b00110110 ;
			12'h00000D04 : data <= 8'b00110110 ;
			12'h00000D05 : data <= 8'b00110110 ;
			12'h00000D06 : data <= 8'b00110110 ;
			12'h00000D07 : data <= 8'b11111111 ;
			12'h00000D08 : data <= 8'b00000000 ;
			12'h00000D09 : data <= 8'b00000000 ;
			12'h00000D0A : data <= 8'b00000000 ;
			12'h00000D0B : data <= 8'b00000000 ;
			12'h00000D0C : data <= 8'b00000000 ;
			12'h00000D0D : data <= 8'b00000000 ;
			12'h00000D0E : data <= 8'b00000000 ;
			12'h00000D0F : data <= 8'b00000000 ;
			12'h00000D10 : data <= 8'b00000000 ;
			12'h00000D11 : data <= 8'b00000000 ;
			12'h00000D12 : data <= 8'b00000000 ;
			12'h00000D13 : data <= 8'b00000000 ;
			12'h00000D14 : data <= 8'b00000000 ;
			12'h00000D15 : data <= 8'b11111111 ;
			12'h00000D16 : data <= 8'b00000000 ;
			12'h00000D17 : data <= 8'b11111111 ;
			12'h00000D18 : data <= 8'b00011000 ;
			12'h00000D19 : data <= 8'b00011000 ;
			12'h00000D1A : data <= 8'b00011000 ;
			12'h00000D1B : data <= 8'b00011000 ;
			12'h00000D1C : data <= 8'b00011000 ;
			12'h00000D1D : data <= 8'b00011000 ;
			12'h00000D1E : data <= 8'b00011000 ;
			12'h00000D1F : data <= 8'b00011000 ;
			12'h00000D20 : data <= 8'b00000000 ;
			12'h00000D21 : data <= 8'b00000000 ;
			12'h00000D22 : data <= 8'b00000000 ;
			12'h00000D23 : data <= 8'b00000000 ;
			12'h00000D24 : data <= 8'b00000000 ;
			12'h00000D25 : data <= 8'b00000000 ;
			12'h00000D26 : data <= 8'b00000000 ;
			12'h00000D27 : data <= 8'b11111111 ;
			12'h00000D28 : data <= 8'b00110110 ;
			12'h00000D29 : data <= 8'b00110110 ;
			12'h00000D2A : data <= 8'b00110110 ;
			12'h00000D2B : data <= 8'b00110110 ;
			12'h00000D2C : data <= 8'b00110110 ;
			12'h00000D2D : data <= 8'b00110110 ;
			12'h00000D2E : data <= 8'b00110110 ;
			12'h00000D2F : data <= 8'b00110110 ;
			12'h00000D30 : data <= 8'b00110110 ;
			12'h00000D31 : data <= 8'b00110110 ;
			12'h00000D32 : data <= 8'b00110110 ;
			12'h00000D33 : data <= 8'b00110110 ;
			12'h00000D34 : data <= 8'b00110110 ;
			12'h00000D35 : data <= 8'b00110110 ;
			12'h00000D36 : data <= 8'b00110110 ;
			12'h00000D37 : data <= 8'b00111111 ;
			12'h00000D38 : data <= 8'b00000000 ;
			12'h00000D39 : data <= 8'b00000000 ;
			12'h00000D3A : data <= 8'b00000000 ;
			12'h00000D3B : data <= 8'b00000000 ;
			12'h00000D3C : data <= 8'b00000000 ;
			12'h00000D3D : data <= 8'b00000000 ;
			12'h00000D3E : data <= 8'b00000000 ;
			12'h00000D3F : data <= 8'b00000000 ;
			12'h00000D40 : data <= 8'b00011000 ;
			12'h00000D41 : data <= 8'b00011000 ;
			12'h00000D42 : data <= 8'b00011000 ;
			12'h00000D43 : data <= 8'b00011000 ;
			12'h00000D44 : data <= 8'b00011000 ;
			12'h00000D45 : data <= 8'b00011111 ;
			12'h00000D46 : data <= 8'b00011000 ;
			12'h00000D47 : data <= 8'b00011111 ;
			12'h00000D48 : data <= 8'b00000000 ;
			12'h00000D49 : data <= 8'b00000000 ;
			12'h00000D4A : data <= 8'b00000000 ;
			12'h00000D4B : data <= 8'b00000000 ;
			12'h00000D4C : data <= 8'b00000000 ;
			12'h00000D4D : data <= 8'b00000000 ;
			12'h00000D4E : data <= 8'b00000000 ;
			12'h00000D4F : data <= 8'b00000000 ;
			12'h00000D50 : data <= 8'b00000000 ;
			12'h00000D51 : data <= 8'b00000000 ;
			12'h00000D52 : data <= 8'b00000000 ;
			12'h00000D53 : data <= 8'b00000000 ;
			12'h00000D54 : data <= 8'b00000000 ;
			12'h00000D55 : data <= 8'b00011111 ;
			12'h00000D56 : data <= 8'b00011000 ;
			12'h00000D57 : data <= 8'b00011111 ;
			12'h00000D58 : data <= 8'b00011000 ;
			12'h00000D59 : data <= 8'b00011000 ;
			12'h00000D5A : data <= 8'b00011000 ;
			12'h00000D5B : data <= 8'b00011000 ;
			12'h00000D5C : data <= 8'b00011000 ;
			12'h00000D5D : data <= 8'b00011000 ;
			12'h00000D5E : data <= 8'b00011000 ;
			12'h00000D5F : data <= 8'b00011000 ;
			12'h00000D60 : data <= 8'b00000000 ;
			12'h00000D61 : data <= 8'b00000000 ;
			12'h00000D62 : data <= 8'b00000000 ;
			12'h00000D63 : data <= 8'b00000000 ;
			12'h00000D64 : data <= 8'b00000000 ;
			12'h00000D65 : data <= 8'b00000000 ;
			12'h00000D66 : data <= 8'b00000000 ;
			12'h00000D67 : data <= 8'b00111111 ;
			12'h00000D68 : data <= 8'b00110110 ;
			12'h00000D69 : data <= 8'b00110110 ;
			12'h00000D6A : data <= 8'b00110110 ;
			12'h00000D6B : data <= 8'b00110110 ;
			12'h00000D6C : data <= 8'b00110110 ;
			12'h00000D6D : data <= 8'b00110110 ;
			12'h00000D6E : data <= 8'b00110110 ;
			12'h00000D6F : data <= 8'b00110110 ;
			12'h00000D70 : data <= 8'b00110110 ;
			12'h00000D71 : data <= 8'b00110110 ;
			12'h00000D72 : data <= 8'b00110110 ;
			12'h00000D73 : data <= 8'b00110110 ;
			12'h00000D74 : data <= 8'b00110110 ;
			12'h00000D75 : data <= 8'b00110110 ;
			12'h00000D76 : data <= 8'b00110110 ;
			12'h00000D77 : data <= 8'b11111111 ;
			12'h00000D78 : data <= 8'b00110110 ;
			12'h00000D79 : data <= 8'b00110110 ;
			12'h00000D7A : data <= 8'b00110110 ;
			12'h00000D7B : data <= 8'b00110110 ;
			12'h00000D7C : data <= 8'b00110110 ;
			12'h00000D7D : data <= 8'b00110110 ;
			12'h00000D7E : data <= 8'b00110110 ;
			12'h00000D7F : data <= 8'b00110110 ;
			12'h00000D80 : data <= 8'b00011000 ;
			12'h00000D81 : data <= 8'b00011000 ;
			12'h00000D82 : data <= 8'b00011000 ;
			12'h00000D83 : data <= 8'b00011000 ;
			12'h00000D84 : data <= 8'b00011000 ;
			12'h00000D85 : data <= 8'b11111111 ;
			12'h00000D86 : data <= 8'b00011000 ;
			12'h00000D87 : data <= 8'b11111111 ;
			12'h00000D88 : data <= 8'b00011000 ;
			12'h00000D89 : data <= 8'b00011000 ;
			12'h00000D8A : data <= 8'b00011000 ;
			12'h00000D8B : data <= 8'b00011000 ;
			12'h00000D8C : data <= 8'b00011000 ;
			12'h00000D8D : data <= 8'b00011000 ;
			12'h00000D8E : data <= 8'b00011000 ;
			12'h00000D8F : data <= 8'b00011000 ;
			12'h00000D90 : data <= 8'b00011000 ;
			12'h00000D91 : data <= 8'b00011000 ;
			12'h00000D92 : data <= 8'b00011000 ;
			12'h00000D93 : data <= 8'b00011000 ;
			12'h00000D94 : data <= 8'b00011000 ;
			12'h00000D95 : data <= 8'b00011000 ;
			12'h00000D96 : data <= 8'b00011000 ;
			12'h00000D97 : data <= 8'b11111000 ;
			12'h00000D98 : data <= 8'b00000000 ;
			12'h00000D99 : data <= 8'b00000000 ;
			12'h00000D9A : data <= 8'b00000000 ;
			12'h00000D9B : data <= 8'b00000000 ;
			12'h00000D9C : data <= 8'b00000000 ;
			12'h00000D9D : data <= 8'b00000000 ;
			12'h00000D9E : data <= 8'b00000000 ;
			12'h00000D9F : data <= 8'b00000000 ;
			12'h00000DA0 : data <= 8'b00000000 ;
			12'h00000DA1 : data <= 8'b00000000 ;
			12'h00000DA2 : data <= 8'b00000000 ;
			12'h00000DA3 : data <= 8'b00000000 ;
			12'h00000DA4 : data <= 8'b00000000 ;
			12'h00000DA5 : data <= 8'b00000000 ;
			12'h00000DA6 : data <= 8'b00000000 ;
			12'h00000DA7 : data <= 8'b00011111 ;
			12'h00000DA8 : data <= 8'b00011000 ;
			12'h00000DA9 : data <= 8'b00011000 ;
			12'h00000DAA : data <= 8'b00011000 ;
			12'h00000DAB : data <= 8'b00011000 ;
			12'h00000DAC : data <= 8'b00011000 ;
			12'h00000DAD : data <= 8'b00011000 ;
			12'h00000DAE : data <= 8'b00011000 ;
			12'h00000DAF : data <= 8'b00011000 ;
			12'h00000DB0 : data <= 8'b11111111 ;
			12'h00000DB1 : data <= 8'b11111111 ;
			12'h00000DB2 : data <= 8'b11111111 ;
			12'h00000DB3 : data <= 8'b11111111 ;
			12'h00000DB4 : data <= 8'b11111111 ;
			12'h00000DB5 : data <= 8'b11111111 ;
			12'h00000DB6 : data <= 8'b11111111 ;
			12'h00000DB7 : data <= 8'b11111111 ;
			12'h00000DB8 : data <= 8'b11111111 ;
			12'h00000DB9 : data <= 8'b11111111 ;
			12'h00000DBA : data <= 8'b11111111 ;
			12'h00000DBB : data <= 8'b11111111 ;
			12'h00000DBC : data <= 8'b11111111 ;
			12'h00000DBD : data <= 8'b11111111 ;
			12'h00000DBE : data <= 8'b11111111 ;
			12'h00000DBF : data <= 8'b11111111 ;
			12'h00000DC0 : data <= 8'b00000000 ;
			12'h00000DC1 : data <= 8'b00000000 ;
			12'h00000DC2 : data <= 8'b00000000 ;
			12'h00000DC3 : data <= 8'b00000000 ;
			12'h00000DC4 : data <= 8'b00000000 ;
			12'h00000DC5 : data <= 8'b00000000 ;
			12'h00000DC6 : data <= 8'b00000000 ;
			12'h00000DC7 : data <= 8'b11111111 ;
			12'h00000DC8 : data <= 8'b11111111 ;
			12'h00000DC9 : data <= 8'b11111111 ;
			12'h00000DCA : data <= 8'b11111111 ;
			12'h00000DCB : data <= 8'b11111111 ;
			12'h00000DCC : data <= 8'b11111111 ;
			12'h00000DCD : data <= 8'b11111111 ;
			12'h00000DCE : data <= 8'b11111111 ;
			12'h00000DCF : data <= 8'b11111111 ;
			12'h00000DD0 : data <= 8'b11110000 ;
			12'h00000DD1 : data <= 8'b11110000 ;
			12'h00000DD2 : data <= 8'b11110000 ;
			12'h00000DD3 : data <= 8'b11110000 ;
			12'h00000DD4 : data <= 8'b11110000 ;
			12'h00000DD5 : data <= 8'b11110000 ;
			12'h00000DD6 : data <= 8'b11110000 ;
			12'h00000DD7 : data <= 8'b11110000 ;
			12'h00000DD8 : data <= 8'b11110000 ;
			12'h00000DD9 : data <= 8'b11110000 ;
			12'h00000DDA : data <= 8'b11110000 ;
			12'h00000DDB : data <= 8'b11110000 ;
			12'h00000DDC : data <= 8'b11110000 ;
			12'h00000DDD : data <= 8'b11110000 ;
			12'h00000DDE : data <= 8'b11110000 ;
			12'h00000DDF : data <= 8'b11110000 ;
			12'h00000DE0 : data <= 8'b00001111 ;
			12'h00000DE1 : data <= 8'b00001111 ;
			12'h00000DE2 : data <= 8'b00001111 ;
			12'h00000DE3 : data <= 8'b00001111 ;
			12'h00000DE4 : data <= 8'b00001111 ;
			12'h00000DE5 : data <= 8'b00001111 ;
			12'h00000DE6 : data <= 8'b00001111 ;
			12'h00000DE7 : data <= 8'b00001111 ;
			12'h00000DE8 : data <= 8'b00001111 ;
			12'h00000DE9 : data <= 8'b00001111 ;
			12'h00000DEA : data <= 8'b00001111 ;
			12'h00000DEB : data <= 8'b00001111 ;
			12'h00000DEC : data <= 8'b00001111 ;
			12'h00000DED : data <= 8'b00001111 ;
			12'h00000DEE : data <= 8'b00001111 ;
			12'h00000DEF : data <= 8'b00001111 ;
			12'h00000DF0 : data <= 8'b11111111 ;
			12'h00000DF1 : data <= 8'b11111111 ;
			12'h00000DF2 : data <= 8'b11111111 ;
			12'h00000DF3 : data <= 8'b11111111 ;
			12'h00000DF4 : data <= 8'b11111111 ;
			12'h00000DF5 : data <= 8'b11111111 ;
			12'h00000DF6 : data <= 8'b11111111 ;
			12'h00000DF7 : data <= 8'b00000000 ;
			12'h00000DF8 : data <= 8'b00000000 ;
			12'h00000DF9 : data <= 8'b00000000 ;
			12'h00000DFA : data <= 8'b00000000 ;
			12'h00000DFB : data <= 8'b00000000 ;
			12'h00000DFC : data <= 8'b00000000 ;
			12'h00000DFD : data <= 8'b00000000 ;
			12'h00000DFE : data <= 8'b00000000 ;
			12'h00000DFF : data <= 8'b00000000 ;
			12'h00000E00 : data <= 8'b00000000 ;
			12'h00000E01 : data <= 8'b00000000 ;
			12'h00000E02 : data <= 8'b00000000 ;
			12'h00000E03 : data <= 8'b00000000 ;
			12'h00000E04 : data <= 8'b00000000 ;
			12'h00000E05 : data <= 8'b01110110 ;
			12'h00000E06 : data <= 8'b11011100 ;
			12'h00000E07 : data <= 8'b11011000 ;
			12'h00000E08 : data <= 8'b11011000 ;
			12'h00000E09 : data <= 8'b11011000 ;
			12'h00000E0A : data <= 8'b11011100 ;
			12'h00000E0B : data <= 8'b01110110 ;
			12'h00000E0C : data <= 8'b00000000 ;
			12'h00000E0D : data <= 8'b00000000 ;
			12'h00000E0E : data <= 8'b00000000 ;
			12'h00000E0F : data <= 8'b00000000 ;
			12'h00000E10 : data <= 8'b00000000 ;
			12'h00000E11 : data <= 8'b00000000 ;
			12'h00000E12 : data <= 8'b01111000 ;
			12'h00000E13 : data <= 8'b11001100 ;
			12'h00000E14 : data <= 8'b11001100 ;
			12'h00000E15 : data <= 8'b11001100 ;
			12'h00000E16 : data <= 8'b11011000 ;
			12'h00000E17 : data <= 8'b11001100 ;
			12'h00000E18 : data <= 8'b11000110 ;
			12'h00000E19 : data <= 8'b11000110 ;
			12'h00000E1A : data <= 8'b11000110 ;
			12'h00000E1B : data <= 8'b11001100 ;
			12'h00000E1C : data <= 8'b00000000 ;
			12'h00000E1D : data <= 8'b00000000 ;
			12'h00000E1E : data <= 8'b00000000 ;
			12'h00000E1F : data <= 8'b00000000 ;
			12'h00000E20 : data <= 8'b00000000 ;
			12'h00000E21 : data <= 8'b00000000 ;
			12'h00000E22 : data <= 8'b11111110 ;
			12'h00000E23 : data <= 8'b11000110 ;
			12'h00000E24 : data <= 8'b11000110 ;
			12'h00000E25 : data <= 8'b11000000 ;
			12'h00000E26 : data <= 8'b11000000 ;
			12'h00000E27 : data <= 8'b11000000 ;
			12'h00000E28 : data <= 8'b11000000 ;
			12'h00000E29 : data <= 8'b11000000 ;
			12'h00000E2A : data <= 8'b11000000 ;
			12'h00000E2B : data <= 8'b11000000 ;
			12'h00000E2C : data <= 8'b00000000 ;
			12'h00000E2D : data <= 8'b00000000 ;
			12'h00000E2E : data <= 8'b00000000 ;
			12'h00000E2F : data <= 8'b00000000 ;
			12'h00000E30 : data <= 8'b00000000 ;
			12'h00000E31 : data <= 8'b00000000 ;
			12'h00000E32 : data <= 8'b00000000 ;
			12'h00000E33 : data <= 8'b00000000 ;
			12'h00000E34 : data <= 8'b11111110 ;
			12'h00000E35 : data <= 8'b01101100 ;
			12'h00000E36 : data <= 8'b01101100 ;
			12'h00000E37 : data <= 8'b01101100 ;
			12'h00000E38 : data <= 8'b01101100 ;
			12'h00000E39 : data <= 8'b01101100 ;
			12'h00000E3A : data <= 8'b01101100 ;
			12'h00000E3B : data <= 8'b01101100 ;
			12'h00000E3C : data <= 8'b00000000 ;
			12'h00000E3D : data <= 8'b00000000 ;
			12'h00000E3E : data <= 8'b00000000 ;
			12'h00000E3F : data <= 8'b00000000 ;
			12'h00000E40 : data <= 8'b00000000 ;
			12'h00000E41 : data <= 8'b00000000 ;
			12'h00000E42 : data <= 8'b00000000 ;
			12'h00000E43 : data <= 8'b11111110 ;
			12'h00000E44 : data <= 8'b11000110 ;
			12'h00000E45 : data <= 8'b01100000 ;
			12'h00000E46 : data <= 8'b00110000 ;
			12'h00000E47 : data <= 8'b00011000 ;
			12'h00000E48 : data <= 8'b00110000 ;
			12'h00000E49 : data <= 8'b01100000 ;
			12'h00000E4A : data <= 8'b11000110 ;
			12'h00000E4B : data <= 8'b11111110 ;
			12'h00000E4C : data <= 8'b00000000 ;
			12'h00000E4D : data <= 8'b00000000 ;
			12'h00000E4E : data <= 8'b00000000 ;
			12'h00000E4F : data <= 8'b00000000 ;
			12'h00000E50 : data <= 8'b00000000 ;
			12'h00000E51 : data <= 8'b00000000 ;
			12'h00000E52 : data <= 8'b00000000 ;
			12'h00000E53 : data <= 8'b00000000 ;
			12'h00000E54 : data <= 8'b00000000 ;
			12'h00000E55 : data <= 8'b01111110 ;
			12'h00000E56 : data <= 8'b11011000 ;
			12'h00000E57 : data <= 8'b11011000 ;
			12'h00000E58 : data <= 8'b11011000 ;
			12'h00000E59 : data <= 8'b11011000 ;
			12'h00000E5A : data <= 8'b11011000 ;
			12'h00000E5B : data <= 8'b01110000 ;
			12'h00000E5C : data <= 8'b00000000 ;
			12'h00000E5D : data <= 8'b00000000 ;
			12'h00000E5E : data <= 8'b00000000 ;
			12'h00000E5F : data <= 8'b00000000 ;
			12'h00000E60 : data <= 8'b00000000 ;
			12'h00000E61 : data <= 8'b00000000 ;
			12'h00000E62 : data <= 8'b00000000 ;
			12'h00000E63 : data <= 8'b00000000 ;
			12'h00000E64 : data <= 8'b01100110 ;
			12'h00000E65 : data <= 8'b01100110 ;
			12'h00000E66 : data <= 8'b01100110 ;
			12'h00000E67 : data <= 8'b01100110 ;
			12'h00000E68 : data <= 8'b01100110 ;
			12'h00000E69 : data <= 8'b01111100 ;
			12'h00000E6A : data <= 8'b01100000 ;
			12'h00000E6B : data <= 8'b01100000 ;
			12'h00000E6C : data <= 8'b11000000 ;
			12'h00000E6D : data <= 8'b00000000 ;
			12'h00000E6E : data <= 8'b00000000 ;
			12'h00000E6F : data <= 8'b00000000 ;
			12'h00000E70 : data <= 8'b00000000 ;
			12'h00000E71 : data <= 8'b00000000 ;
			12'h00000E72 : data <= 8'b00000000 ;
			12'h00000E73 : data <= 8'b00000000 ;
			12'h00000E74 : data <= 8'b01110110 ;
			12'h00000E75 : data <= 8'b11011100 ;
			12'h00000E76 : data <= 8'b00011000 ;
			12'h00000E77 : data <= 8'b00011000 ;
			12'h00000E78 : data <= 8'b00011000 ;
			12'h00000E79 : data <= 8'b00011000 ;
			12'h00000E7A : data <= 8'b00011000 ;
			12'h00000E7B : data <= 8'b00011000 ;
			12'h00000E7C : data <= 8'b00000000 ;
			12'h00000E7D : data <= 8'b00000000 ;
			12'h00000E7E : data <= 8'b00000000 ;
			12'h00000E7F : data <= 8'b00000000 ;
			12'h00000E80 : data <= 8'b00000000 ;
			12'h00000E81 : data <= 8'b00000000 ;
			12'h00000E82 : data <= 8'b00000000 ;
			12'h00000E83 : data <= 8'b01111110 ;
			12'h00000E84 : data <= 8'b00011000 ;
			12'h00000E85 : data <= 8'b00111100 ;
			12'h00000E86 : data <= 8'b01100110 ;
			12'h00000E87 : data <= 8'b01100110 ;
			12'h00000E88 : data <= 8'b01100110 ;
			12'h00000E89 : data <= 8'b00111100 ;
			12'h00000E8A : data <= 8'b00011000 ;
			12'h00000E8B : data <= 8'b01111110 ;
			12'h00000E8C : data <= 8'b00000000 ;
			12'h00000E8D : data <= 8'b00000000 ;
			12'h00000E8E : data <= 8'b00000000 ;
			12'h00000E8F : data <= 8'b00000000 ;
			12'h00000E90 : data <= 8'b00000000 ;
			12'h00000E91 : data <= 8'b00000000 ;
			12'h00000E92 : data <= 8'b00000000 ;
			12'h00000E93 : data <= 8'b00111000 ;
			12'h00000E94 : data <= 8'b01101100 ;
			12'h00000E95 : data <= 8'b11000110 ;
			12'h00000E96 : data <= 8'b11000110 ;
			12'h00000E97 : data <= 8'b11111110 ;
			12'h00000E98 : data <= 8'b11000110 ;
			12'h00000E99 : data <= 8'b11000110 ;
			12'h00000E9A : data <= 8'b01101100 ;
			12'h00000E9B : data <= 8'b00111000 ;
			12'h00000E9C : data <= 8'b00000000 ;
			12'h00000E9D : data <= 8'b00000000 ;
			12'h00000E9E : data <= 8'b00000000 ;
			12'h00000E9F : data <= 8'b00000000 ;
			12'h00000EA0 : data <= 8'b00000000 ;
			12'h00000EA1 : data <= 8'b00000000 ;
			12'h00000EA2 : data <= 8'b00111000 ;
			12'h00000EA3 : data <= 8'b01101100 ;
			12'h00000EA4 : data <= 8'b11000110 ;
			12'h00000EA5 : data <= 8'b11000110 ;
			12'h00000EA6 : data <= 8'b11000110 ;
			12'h00000EA7 : data <= 8'b01101100 ;
			12'h00000EA8 : data <= 8'b01101100 ;
			12'h00000EA9 : data <= 8'b01101100 ;
			12'h00000EAA : data <= 8'b01101100 ;
			12'h00000EAB : data <= 8'b11101110 ;
			12'h00000EAC : data <= 8'b00000000 ;
			12'h00000EAD : data <= 8'b00000000 ;
			12'h00000EAE : data <= 8'b00000000 ;
			12'h00000EAF : data <= 8'b00000000 ;
			12'h00000EB0 : data <= 8'b00000000 ;
			12'h00000EB1 : data <= 8'b00000000 ;
			12'h00000EB2 : data <= 8'b00011110 ;
			12'h00000EB3 : data <= 8'b00110000 ;
			12'h00000EB4 : data <= 8'b00011000 ;
			12'h00000EB5 : data <= 8'b00001100 ;
			12'h00000EB6 : data <= 8'b00111110 ;
			12'h00000EB7 : data <= 8'b01100110 ;
			12'h00000EB8 : data <= 8'b01100110 ;
			12'h00000EB9 : data <= 8'b01100110 ;
			12'h00000EBA : data <= 8'b01100110 ;
			12'h00000EBB : data <= 8'b00111100 ;
			12'h00000EBC : data <= 8'b00000000 ;
			12'h00000EBD : data <= 8'b00000000 ;
			12'h00000EBE : data <= 8'b00000000 ;
			12'h00000EBF : data <= 8'b00000000 ;
			12'h00000EC0 : data <= 8'b00000000 ;
			12'h00000EC1 : data <= 8'b00000000 ;
			12'h00000EC2 : data <= 8'b00000000 ;
			12'h00000EC3 : data <= 8'b00000000 ;
			12'h00000EC4 : data <= 8'b00000000 ;
			12'h00000EC5 : data <= 8'b01111110 ;
			12'h00000EC6 : data <= 8'b11011011 ;
			12'h00000EC7 : data <= 8'b11011011 ;
			12'h00000EC8 : data <= 8'b11011011 ;
			12'h00000EC9 : data <= 8'b01111110 ;
			12'h00000ECA : data <= 8'b00000000 ;
			12'h00000ECB : data <= 8'b00000000 ;
			12'h00000ECC : data <= 8'b00000000 ;
			12'h00000ECD : data <= 8'b00000000 ;
			12'h00000ECE : data <= 8'b00000000 ;
			12'h00000ECF : data <= 8'b00000000 ;
			12'h00000ED0 : data <= 8'b00000000 ;
			12'h00000ED1 : data <= 8'b00000000 ;
			12'h00000ED2 : data <= 8'b00000000 ;
			12'h00000ED3 : data <= 8'b00000011 ;
			12'h00000ED4 : data <= 8'b00000110 ;
			12'h00000ED5 : data <= 8'b01111110 ;
			12'h00000ED6 : data <= 8'b11011011 ;
			12'h00000ED7 : data <= 8'b11011011 ;
			12'h00000ED8 : data <= 8'b11110011 ;
			12'h00000ED9 : data <= 8'b01111110 ;
			12'h00000EDA : data <= 8'b01100000 ;
			12'h00000EDB : data <= 8'b11000000 ;
			12'h00000EDC : data <= 8'b00000000 ;
			12'h00000EDD : data <= 8'b00000000 ;
			12'h00000EDE : data <= 8'b00000000 ;
			12'h00000EDF : data <= 8'b00000000 ;
			12'h00000EE0 : data <= 8'b00000000 ;
			12'h00000EE1 : data <= 8'b00000000 ;
			12'h00000EE2 : data <= 8'b00011100 ;
			12'h00000EE3 : data <= 8'b00110000 ;
			12'h00000EE4 : data <= 8'b01100000 ;
			12'h00000EE5 : data <= 8'b01100000 ;
			12'h00000EE6 : data <= 8'b01111100 ;
			12'h00000EE7 : data <= 8'b01100000 ;
			12'h00000EE8 : data <= 8'b01100000 ;
			12'h00000EE9 : data <= 8'b01100000 ;
			12'h00000EEA : data <= 8'b00110000 ;
			12'h00000EEB : data <= 8'b00011100 ;
			12'h00000EEC : data <= 8'b00000000 ;
			12'h00000EED : data <= 8'b00000000 ;
			12'h00000EEE : data <= 8'b00000000 ;
			12'h00000EEF : data <= 8'b00000000 ;
			12'h00000EF0 : data <= 8'b00000000 ;
			12'h00000EF1 : data <= 8'b00000000 ;
			12'h00000EF2 : data <= 8'b00000000 ;
			12'h00000EF3 : data <= 8'b01111100 ;
			12'h00000EF4 : data <= 8'b11000110 ;
			12'h00000EF5 : data <= 8'b11000110 ;
			12'h00000EF6 : data <= 8'b11000110 ;
			12'h00000EF7 : data <= 8'b11000110 ;
			12'h00000EF8 : data <= 8'b11000110 ;
			12'h00000EF9 : data <= 8'b11000110 ;
			12'h00000EFA : data <= 8'b11000110 ;
			12'h00000EFB : data <= 8'b11000110 ;
			12'h00000EFC : data <= 8'b00000000 ;
			12'h00000EFD : data <= 8'b00000000 ;
			12'h00000EFE : data <= 8'b00000000 ;
			12'h00000EFF : data <= 8'b00000000 ;
			12'h00000F00 : data <= 8'b00000000 ;
			12'h00000F01 : data <= 8'b00000000 ;
			12'h00000F02 : data <= 8'b00000000 ;
			12'h00000F03 : data <= 8'b00000000 ;
			12'h00000F04 : data <= 8'b11111110 ;
			12'h00000F05 : data <= 8'b00000000 ;
			12'h00000F06 : data <= 8'b00000000 ;
			12'h00000F07 : data <= 8'b11111110 ;
			12'h00000F08 : data <= 8'b00000000 ;
			12'h00000F09 : data <= 8'b00000000 ;
			12'h00000F0A : data <= 8'b11111110 ;
			12'h00000F0B : data <= 8'b00000000 ;
			12'h00000F0C : data <= 8'b00000000 ;
			12'h00000F0D : data <= 8'b00000000 ;
			12'h00000F0E : data <= 8'b00000000 ;
			12'h00000F0F : data <= 8'b00000000 ;
			12'h00000F10 : data <= 8'b00000000 ;
			12'h00000F11 : data <= 8'b00000000 ;
			12'h00000F12 : data <= 8'b00000000 ;
			12'h00000F13 : data <= 8'b00000000 ;
			12'h00000F14 : data <= 8'b00011000 ;
			12'h00000F15 : data <= 8'b00011000 ;
			12'h00000F16 : data <= 8'b01111110 ;
			12'h00000F17 : data <= 8'b00011000 ;
			12'h00000F18 : data <= 8'b00011000 ;
			12'h00000F19 : data <= 8'b00000000 ;
			12'h00000F1A : data <= 8'b00000000 ;
			12'h00000F1B : data <= 8'b11111111 ;
			12'h00000F1C : data <= 8'b00000000 ;
			12'h00000F1D : data <= 8'b00000000 ;
			12'h00000F1E : data <= 8'b00000000 ;
			12'h00000F1F : data <= 8'b00000000 ;
			12'h00000F20 : data <= 8'b00000000 ;
			12'h00000F21 : data <= 8'b00000000 ;
			12'h00000F22 : data <= 8'b00000000 ;
			12'h00000F23 : data <= 8'b00110000 ;
			12'h00000F24 : data <= 8'b00011000 ;
			12'h00000F25 : data <= 8'b00001100 ;
			12'h00000F26 : data <= 8'b00000110 ;
			12'h00000F27 : data <= 8'b00001100 ;
			12'h00000F28 : data <= 8'b00011000 ;
			12'h00000F29 : data <= 8'b00110000 ;
			12'h00000F2A : data <= 8'b00000000 ;
			12'h00000F2B : data <= 8'b01111110 ;
			12'h00000F2C : data <= 8'b00000000 ;
			12'h00000F2D : data <= 8'b00000000 ;
			12'h00000F2E : data <= 8'b00000000 ;
			12'h00000F2F : data <= 8'b00000000 ;
			12'h00000F30 : data <= 8'b00000000 ;
			12'h00000F31 : data <= 8'b00000000 ;
			12'h00000F32 : data <= 8'b00000000 ;
			12'h00000F33 : data <= 8'b00001100 ;
			12'h00000F34 : data <= 8'b00011000 ;
			12'h00000F35 : data <= 8'b00110000 ;
			12'h00000F36 : data <= 8'b01100000 ;
			12'h00000F37 : data <= 8'b00110000 ;
			12'h00000F38 : data <= 8'b00011000 ;
			12'h00000F39 : data <= 8'b00001100 ;
			12'h00000F3A : data <= 8'b00000000 ;
			12'h00000F3B : data <= 8'b01111110 ;
			12'h00000F3C : data <= 8'b00000000 ;
			12'h00000F3D : data <= 8'b00000000 ;
			12'h00000F3E : data <= 8'b00000000 ;
			12'h00000F3F : data <= 8'b00000000 ;
			12'h00000F40 : data <= 8'b00000000 ;
			12'h00000F41 : data <= 8'b00000000 ;
			12'h00000F42 : data <= 8'b00001110 ;
			12'h00000F43 : data <= 8'b00011011 ;
			12'h00000F44 : data <= 8'b00011011 ;
			12'h00000F45 : data <= 8'b00011000 ;
			12'h00000F46 : data <= 8'b00011000 ;
			12'h00000F47 : data <= 8'b00011000 ;
			12'h00000F48 : data <= 8'b00011000 ;
			12'h00000F49 : data <= 8'b00011000 ;
			12'h00000F4A : data <= 8'b00011000 ;
			12'h00000F4B : data <= 8'b00011000 ;
			12'h00000F4C : data <= 8'b00011000 ;
			12'h00000F4D : data <= 8'b00011000 ;
			12'h00000F4E : data <= 8'b00011000 ;
			12'h00000F4F : data <= 8'b00011000 ;
			12'h00000F50 : data <= 8'b00011000 ;
			12'h00000F51 : data <= 8'b00011000 ;
			12'h00000F52 : data <= 8'b00011000 ;
			12'h00000F53 : data <= 8'b00011000 ;
			12'h00000F54 : data <= 8'b00011000 ;
			12'h00000F55 : data <= 8'b00011000 ;
			12'h00000F56 : data <= 8'b00011000 ;
			12'h00000F57 : data <= 8'b00011000 ;
			12'h00000F58 : data <= 8'b11011000 ;
			12'h00000F59 : data <= 8'b11011000 ;
			12'h00000F5A : data <= 8'b11011000 ;
			12'h00000F5B : data <= 8'b01110000 ;
			12'h00000F5C : data <= 8'b00000000 ;
			12'h00000F5D : data <= 8'b00000000 ;
			12'h00000F5E : data <= 8'b00000000 ;
			12'h00000F5F : data <= 8'b00000000 ;
			12'h00000F60 : data <= 8'b00000000 ;
			12'h00000F61 : data <= 8'b00000000 ;
			12'h00000F62 : data <= 8'b00000000 ;
			12'h00000F63 : data <= 8'b00000000 ;
			12'h00000F64 : data <= 8'b00011000 ;
			12'h00000F65 : data <= 8'b00011000 ;
			12'h00000F66 : data <= 8'b00000000 ;
			12'h00000F67 : data <= 8'b01111110 ;
			12'h00000F68 : data <= 8'b00000000 ;
			12'h00000F69 : data <= 8'b00011000 ;
			12'h00000F6A : data <= 8'b00011000 ;
			12'h00000F6B : data <= 8'b00000000 ;
			12'h00000F6C : data <= 8'b00000000 ;
			12'h00000F6D : data <= 8'b00000000 ;
			12'h00000F6E : data <= 8'b00000000 ;
			12'h00000F6F : data <= 8'b00000000 ;
			12'h00000F70 : data <= 8'b00000000 ;
			12'h00000F71 : data <= 8'b00000000 ;
			12'h00000F72 : data <= 8'b00000000 ;
			12'h00000F73 : data <= 8'b00000000 ;
			12'h00000F74 : data <= 8'b00000000 ;
			12'h00000F75 : data <= 8'b01110110 ;
			12'h00000F76 : data <= 8'b11011100 ;
			12'h00000F77 : data <= 8'b00000000 ;
			12'h00000F78 : data <= 8'b01110110 ;
			12'h00000F79 : data <= 8'b11011100 ;
			12'h00000F7A : data <= 8'b00000000 ;
			12'h00000F7B : data <= 8'b00000000 ;
			12'h00000F7C : data <= 8'b00000000 ;
			12'h00000F7D : data <= 8'b00000000 ;
			12'h00000F7E : data <= 8'b00000000 ;
			12'h00000F7F : data <= 8'b00000000 ;
			12'h00000F80 : data <= 8'b00000000 ;
			12'h00000F81 : data <= 8'b00111000 ;
			12'h00000F82 : data <= 8'b01101100 ;
			12'h00000F83 : data <= 8'b01101100 ;
			12'h00000F84 : data <= 8'b00111000 ;
			12'h00000F85 : data <= 8'b00000000 ;
			12'h00000F86 : data <= 8'b00000000 ;
			12'h00000F87 : data <= 8'b00000000 ;
			12'h00000F88 : data <= 8'b00000000 ;
			12'h00000F89 : data <= 8'b00000000 ;
			12'h00000F8A : data <= 8'b00000000 ;
			12'h00000F8B : data <= 8'b00000000 ;
			12'h00000F8C : data <= 8'b00000000 ;
			12'h00000F8D : data <= 8'b00000000 ;
			12'h00000F8E : data <= 8'b00000000 ;
			12'h00000F8F : data <= 8'b00000000 ;
			12'h00000F90 : data <= 8'b00000000 ;
			12'h00000F91 : data <= 8'b00000000 ;
			12'h00000F92 : data <= 8'b00000000 ;
			12'h00000F93 : data <= 8'b00000000 ;
			12'h00000F94 : data <= 8'b00000000 ;
			12'h00000F95 : data <= 8'b00000000 ;
			12'h00000F96 : data <= 8'b00000000 ;
			12'h00000F97 : data <= 8'b00011000 ;
			12'h00000F98 : data <= 8'b00011000 ;
			12'h00000F99 : data <= 8'b00000000 ;
			12'h00000F9A : data <= 8'b00000000 ;
			12'h00000F9B : data <= 8'b00000000 ;
			12'h00000F9C : data <= 8'b00000000 ;
			12'h00000F9D : data <= 8'b00000000 ;
			12'h00000F9E : data <= 8'b00000000 ;
			12'h00000F9F : data <= 8'b00000000 ;
			12'h00000FA0 : data <= 8'b00000000 ;
			12'h00000FA1 : data <= 8'b00000000 ;
			12'h00000FA2 : data <= 8'b00000000 ;
			12'h00000FA3 : data <= 8'b00000000 ;
			12'h00000FA4 : data <= 8'b00000000 ;
			12'h00000FA5 : data <= 8'b00000000 ;
			12'h00000FA6 : data <= 8'b00000000 ;
			12'h00000FA7 : data <= 8'b00000000 ;
			12'h00000FA8 : data <= 8'b00011000 ;
			12'h00000FA9 : data <= 8'b00000000 ;
			12'h00000FAA : data <= 8'b00000000 ;
			12'h00000FAB : data <= 8'b00000000 ;
			12'h00000FAC : data <= 8'b00000000 ;
			12'h00000FAD : data <= 8'b00000000 ;
			12'h00000FAE : data <= 8'b00000000 ;
			12'h00000FAF : data <= 8'b00000000 ;
			12'h00000FB0 : data <= 8'b00000000 ;
			12'h00000FB1 : data <= 8'b00001111 ;
			12'h00000FB2 : data <= 8'b00001100 ;
			12'h00000FB3 : data <= 8'b00001100 ;
			12'h00000FB4 : data <= 8'b00001100 ;
			12'h00000FB5 : data <= 8'b00001100 ;
			12'h00000FB6 : data <= 8'b00001100 ;
			12'h00000FB7 : data <= 8'b11101100 ;
			12'h00000FB8 : data <= 8'b01101100 ;
			12'h00000FB9 : data <= 8'b01101100 ;
			12'h00000FBA : data <= 8'b00111100 ;
			12'h00000FBB : data <= 8'b00011100 ;
			12'h00000FBC : data <= 8'b00000000 ;
			12'h00000FBD : data <= 8'b00000000 ;
			12'h00000FBE : data <= 8'b00000000 ;
			12'h00000FBF : data <= 8'b00000000 ;
			12'h00000FC0 : data <= 8'b00000000 ;
			12'h00000FC1 : data <= 8'b11011000 ;
			12'h00000FC2 : data <= 8'b01101100 ;
			12'h00000FC3 : data <= 8'b01101100 ;
			12'h00000FC4 : data <= 8'b01101100 ;
			12'h00000FC5 : data <= 8'b01101100 ;
			12'h00000FC6 : data <= 8'b01101100 ;
			12'h00000FC7 : data <= 8'b00000000 ;
			12'h00000FC8 : data <= 8'b00000000 ;
			12'h00000FC9 : data <= 8'b00000000 ;
			12'h00000FCA : data <= 8'b00000000 ;
			12'h00000FCB : data <= 8'b00000000 ;
			12'h00000FCC : data <= 8'b00000000 ;
			12'h00000FCD : data <= 8'b00000000 ;
			12'h00000FCE : data <= 8'b00000000 ;
			12'h00000FCF : data <= 8'b00000000 ;
			12'h00000FD0 : data <= 8'b00000000 ;
			12'h00000FD1 : data <= 8'b01110000 ;
			12'h00000FD2 : data <= 8'b11011000 ;
			12'h00000FD3 : data <= 8'b00110000 ;
			12'h00000FD4 : data <= 8'b01100000 ;
			12'h00000FD5 : data <= 8'b11001000 ;
			12'h00000FD6 : data <= 8'b11111000 ;
			12'h00000FD7 : data <= 8'b00000000 ;
			12'h00000FD8 : data <= 8'b00000000 ;
			12'h00000FD9 : data <= 8'b00000000 ;
			12'h00000FDA : data <= 8'b00000000 ;
			12'h00000FDB : data <= 8'b00000000 ;
			12'h00000FDC : data <= 8'b00000000 ;
			12'h00000FDD : data <= 8'b00000000 ;
			12'h00000FDE : data <= 8'b00000000 ;
			12'h00000FDF : data <= 8'b00000000 ;
			12'h00000FE0 : data <= 8'b00000000 ;
			12'h00000FE1 : data <= 8'b00000000 ;
			12'h00000FE2 : data <= 8'b00000000 ;
			12'h00000FE3 : data <= 8'b00000000 ;
			12'h00000FE4 : data <= 8'b01111100 ;
			12'h00000FE5 : data <= 8'b01111100 ;
			12'h00000FE6 : data <= 8'b01111100 ;
			12'h00000FE7 : data <= 8'b01111100 ;
			12'h00000FE8 : data <= 8'b01111100 ;
			12'h00000FE9 : data <= 8'b01111100 ;
			12'h00000FEA : data <= 8'b01111100 ;
			12'h00000FEB : data <= 8'b00000000 ;
			12'h00000FEC : data <= 8'b00000000 ;
			12'h00000FED : data <= 8'b00000000 ;
			12'h00000FEE : data <= 8'b00000000 ;
			12'h00000FEF : data <= 8'b00000000 ;
			12'h00000FF0 : data <= 8'b00000000 ;
			12'h00000FF1 : data <= 8'b00000000 ;
			12'h00000FF2 : data <= 8'b00000000 ;
			12'h00000FF3 : data <= 8'b00000000 ;
			12'h00000FF4 : data <= 8'b00000000 ;
			12'h00000FF5 : data <= 8'b00000000 ;
			12'h00000FF6 : data <= 8'b00000000 ;
			12'h00000FF7 : data <= 8'b00000000 ;
			12'h00000FF8 : data <= 8'b00000000 ;
			12'h00000FF9 : data <= 8'b00000000 ;
			12'h00000FFA : data <= 8'b00000000 ;
			12'h00000FFB : data <= 8'b00000000 ;
			12'h00000FFC : data <= 8'b00000000 ;
			12'h00000FFD : data <= 8'b00000000 ;
			12'h00000FFE : data <= 8'b00000000 ;
			12'h00000FFF : data <= 8'b00000000 ;
		endcase
	end
endmodule